// Generated from: 20251204-054922_binTestAcc8709_seed749733_epochs30_2x8000_b256_lr75_interconnect.npz

module net (
    input  wire [767:0] in,
    output wire [7999:0] out,
    output wire [5109:0] categories
);
    wire [7999:0] layer_0;

    // Layer 0 ============================================================
    assign layer_0[0] = in[107] | in[113]; 
    assign layer_0[1] = in[358]; 
    assign layer_0[2] = ~in[636] | (in[636] & in[118]); 
    assign layer_0[3] = in[43] ^ in[441]; 
    assign layer_0[4] = ~(in[742] & in[373]); 
    assign layer_0[5] = ~in[552] | (in[44] & in[552]); 
    assign layer_0[6] = in[275] | in[676]; 
    assign layer_0[7] = in[744] | in[760]; 
    assign layer_0[8] = 1'b0; 
    assign layer_0[9] = in[505] | in[586]; 
    assign layer_0[10] = ~in[726] | (in[726] & in[522]); 
    assign layer_0[11] = ~(in[4] ^ in[264]); 
    assign layer_0[12] = in[23] & ~in[518]; 
    assign layer_0[13] = in[310] | in[302]; 
    assign layer_0[14] = ~in[310]; 
    assign layer_0[15] = in[499] & in[296]; 
    assign layer_0[16] = in[330] & in[450]; 
    assign layer_0[17] = in[436] ^ in[58]; 
    assign layer_0[18] = ~in[307]; 
    assign layer_0[19] = in[120] & in[313]; 
    assign layer_0[20] = ~in[418] | (in[418] & in[341]); 
    assign layer_0[21] = 1'b0; 
    assign layer_0[22] = in[260] & in[325]; 
    assign layer_0[23] = in[4] ^ in[244]; 
    assign layer_0[24] = ~(in[43] & in[298]); 
    assign layer_0[25] = in[378]; 
    assign layer_0[26] = in[338] ^ in[94]; 
    assign layer_0[27] = in[569] & ~in[491]; 
    assign layer_0[28] = ~(in[551] & in[535]); 
    assign layer_0[29] = ~(in[596] & in[310]); 
    assign layer_0[30] = in[192] ^ in[757]; 
    assign layer_0[31] = in[612]; 
    assign layer_0[32] = in[197] & ~in[676]; 
    assign layer_0[33] = ~(in[597] ^ in[228]); 
    assign layer_0[34] = in[392]; 
    assign layer_0[35] = in[360]; 
    assign layer_0[36] = ~(in[117] & in[293]); 
    assign layer_0[37] = ~in[343]; 
    assign layer_0[38] = in[555]; 
    assign layer_0[39] = in[347] ^ in[633]; 
    assign layer_0[40] = ~(in[109] ^ in[712]); 
    assign layer_0[41] = ~in[179] | (in[525] & in[179]); 
    assign layer_0[42] = ~(in[261] ^ in[680]); 
    assign layer_0[43] = in[501] ^ in[243]; 
    assign layer_0[44] = in[202] | in[638]; 
    assign layer_0[45] = ~(in[331] ^ in[618]); 
    assign layer_0[46] = in[383] | in[206]; 
    assign layer_0[47] = ~in[436] | (in[436] & in[263]); 
    assign layer_0[48] = ~(in[654] ^ in[713]); 
    assign layer_0[49] = ~in[362]; 
    assign layer_0[50] = ~in[618]; 
    assign layer_0[51] = in[660]; 
    assign layer_0[52] = in[725] | in[636]; 
    assign layer_0[53] = in[674] ^ in[662]; 
    assign layer_0[54] = ~(in[363] & in[133]); 
    assign layer_0[55] = in[646] ^ in[601]; 
    assign layer_0[56] = ~(in[284] & in[505]); 
    assign layer_0[57] = in[449] | in[334]; 
    assign layer_0[58] = in[675]; 
    assign layer_0[59] = in[599] ^ in[697]; 
    assign layer_0[60] = ~(in[411] & in[211]); 
    assign layer_0[61] = ~in[378]; 
    assign layer_0[62] = in[293] & ~in[397]; 
    assign layer_0[63] = ~(in[79] ^ in[501]); 
    assign layer_0[64] = ~(in[654] ^ in[717]); 
    assign layer_0[65] = ~in[409] | (in[409] & in[591]); 
    assign layer_0[66] = ~(in[477] | in[368]); 
    assign layer_0[67] = ~(in[541] | in[71]); 
    assign layer_0[68] = in[380]; 
    assign layer_0[69] = in[716]; 
    assign layer_0[70] = in[635]; 
    assign layer_0[71] = in[39] ^ in[267]; 
    assign layer_0[72] = ~(in[634] ^ in[667]); 
    assign layer_0[73] = ~in[331]; 
    assign layer_0[74] = in[100] & ~in[115]; 
    assign layer_0[75] = in[216] & ~in[28]; 
    assign layer_0[76] = ~in[407]; 
    assign layer_0[77] = in[321] | in[297]; 
    assign layer_0[78] = in[623]; 
    assign layer_0[79] = ~(in[611] & in[106]); 
    assign layer_0[80] = ~in[393]; 
    assign layer_0[81] = ~(in[702] ^ in[359]); 
    assign layer_0[82] = ~in[385]; 
    assign layer_0[83] = ~in[452] | (in[452] & in[256]); 
    assign layer_0[84] = ~in[580] | (in[580] & in[699]); 
    assign layer_0[85] = in[52] ^ in[371]; 
    assign layer_0[86] = ~(in[666] & in[643]); 
    assign layer_0[87] = in[400] ^ in[526]; 
    assign layer_0[88] = ~(in[601] | in[298]); 
    assign layer_0[89] = ~in[713]; 
    assign layer_0[90] = 1'b0; 
    assign layer_0[91] = ~(in[509] ^ in[341]); 
    assign layer_0[92] = in[508]; 
    assign layer_0[93] = in[35] & ~in[675]; 
    assign layer_0[94] = ~(in[601] | in[114]); 
    assign layer_0[95] = ~(in[759] ^ in[245]); 
    assign layer_0[96] = ~(in[708] | in[644]); 
    assign layer_0[97] = in[630]; 
    assign layer_0[98] = in[282] ^ in[443]; 
    assign layer_0[99] = ~(in[601] ^ in[3]); 
    assign layer_0[100] = ~in[711] | (in[80] & in[711]); 
    assign layer_0[101] = in[654] & ~in[316]; 
    assign layer_0[102] = in[365] & ~in[222]; 
    assign layer_0[103] = in[669] | in[502]; 
    assign layer_0[104] = in[519] ^ in[276]; 
    assign layer_0[105] = ~(in[173] | in[287]); 
    assign layer_0[106] = ~(in[558] | in[412]); 
    assign layer_0[107] = in[377] | in[304]; 
    assign layer_0[108] = in[71]; 
    assign layer_0[109] = ~(in[382] ^ in[317]); 
    assign layer_0[110] = ~in[619] | (in[500] & in[619]); 
    assign layer_0[111] = in[534] & ~in[275]; 
    assign layer_0[112] = in[273] ^ in[314]; 
    assign layer_0[113] = ~(in[649] | in[47]); 
    assign layer_0[114] = ~in[442]; 
    assign layer_0[115] = ~(in[236] ^ in[128]); 
    assign layer_0[116] = in[223] & ~in[304]; 
    assign layer_0[117] = ~(in[567] ^ in[674]); 
    assign layer_0[118] = ~(in[182] | in[624]); 
    assign layer_0[119] = ~(in[706] ^ in[757]); 
    assign layer_0[120] = ~(in[699] ^ in[676]); 
    assign layer_0[121] = ~(in[221] & in[501]); 
    assign layer_0[122] = in[293]; 
    assign layer_0[123] = ~(in[19] | in[660]); 
    assign layer_0[124] = in[425]; 
    assign layer_0[125] = 1'b1; 
    assign layer_0[126] = ~in[482]; 
    assign layer_0[127] = in[284]; 
    assign layer_0[128] = in[27] & in[56]; 
    assign layer_0[129] = ~(in[759] ^ in[347]); 
    assign layer_0[130] = 1'b1; 
    assign layer_0[131] = in[600] & ~in[167]; 
    assign layer_0[132] = in[400] | in[267]; 
    assign layer_0[133] = ~(in[350] ^ in[568]); 
    assign layer_0[134] = ~(in[760] ^ in[698]); 
    assign layer_0[135] = in[151]; 
    assign layer_0[136] = ~(in[379] | in[346]); 
    assign layer_0[137] = in[195] & in[227]; 
    assign layer_0[138] = ~in[586]; 
    assign layer_0[139] = ~in[282]; 
    assign layer_0[140] = in[702]; 
    assign layer_0[141] = ~(in[603] | in[534]); 
    assign layer_0[142] = ~in[124] | (in[124] & in[628]); 
    assign layer_0[143] = ~in[352] | (in[352] & in[645]); 
    assign layer_0[144] = ~(in[435] ^ in[618]); 
    assign layer_0[145] = ~(in[465] ^ in[449]); 
    assign layer_0[146] = ~(in[111] ^ in[56]); 
    assign layer_0[147] = ~(in[398] ^ in[742]); 
    assign layer_0[148] = ~in[408] | (in[408] & in[762]); 
    assign layer_0[149] = in[266] & ~in[259]; 
    assign layer_0[150] = ~(in[412] ^ in[507]); 
    assign layer_0[151] = ~(in[67] & in[724]); 
    assign layer_0[152] = in[229] & in[584]; 
    assign layer_0[153] = in[129] & in[632]; 
    assign layer_0[154] = in[680] ^ in[341]; 
    assign layer_0[155] = ~(in[242] | in[367]); 
    assign layer_0[156] = ~in[470] | (in[470] & in[499]); 
    assign layer_0[157] = in[449] & ~in[224]; 
    assign layer_0[158] = in[500]; 
    assign layer_0[159] = in[251] ^ in[485]; 
    assign layer_0[160] = in[534] & ~in[539]; 
    assign layer_0[161] = ~(in[580] ^ in[374]); 
    assign layer_0[162] = ~(in[177] ^ in[233]); 
    assign layer_0[163] = ~(in[458] ^ in[580]); 
    assign layer_0[164] = in[483]; 
    assign layer_0[165] = in[450] & ~in[668]; 
    assign layer_0[166] = in[232]; 
    assign layer_0[167] = in[565]; 
    assign layer_0[168] = ~(in[253] & in[695]); 
    assign layer_0[169] = in[500] ^ in[309]; 
    assign layer_0[170] = in[346] & ~in[268]; 
    assign layer_0[171] = 1'b0; 
    assign layer_0[172] = ~(in[618] ^ in[19]); 
    assign layer_0[173] = ~(in[600] & in[475]); 
    assign layer_0[174] = ~in[618]; 
    assign layer_0[175] = in[160] & in[336]; 
    assign layer_0[176] = ~(in[280] ^ in[66]); 
    assign layer_0[177] = in[314] & in[564]; 
    assign layer_0[178] = in[450] ^ in[369]; 
    assign layer_0[179] = ~in[482]; 
    assign layer_0[180] = ~(in[488] & in[109]); 
    assign layer_0[181] = in[7] & in[396]; 
    assign layer_0[182] = in[311] & ~in[324]; 
    assign layer_0[183] = ~in[649]; 
    assign layer_0[184] = in[726] ^ in[600]; 
    assign layer_0[185] = in[493] ^ in[250]; 
    assign layer_0[186] = in[603] & in[421]; 
    assign layer_0[187] = ~in[264] | (in[264] & in[323]); 
    assign layer_0[188] = in[113]; 
    assign layer_0[189] = ~(in[690] ^ in[356]); 
    assign layer_0[190] = ~(in[681] ^ in[550]); 
    assign layer_0[191] = in[346] ^ in[488]; 
    assign layer_0[192] = ~(in[494] ^ in[54]); 
    assign layer_0[193] = ~(in[264] ^ in[18]); 
    assign layer_0[194] = in[284]; 
    assign layer_0[195] = ~(in[268] & in[449]); 
    assign layer_0[196] = ~(in[600] ^ in[28]); 
    assign layer_0[197] = in[127]; 
    assign layer_0[198] = in[446] ^ in[566]; 
    assign layer_0[199] = ~in[727]; 
    assign layer_0[200] = in[399] & ~in[311]; 
    assign layer_0[201] = in[725] ^ in[173]; 
    assign layer_0[202] = ~(in[645] | in[724]); 
    assign layer_0[203] = in[622]; 
    assign layer_0[204] = in[536] & ~in[503]; 
    assign layer_0[205] = ~(in[651] ^ in[44]); 
    assign layer_0[206] = ~(in[371] | in[348]); 
    assign layer_0[207] = in[11] & ~in[605]; 
    assign layer_0[208] = in[568] & ~in[763]; 
    assign layer_0[209] = ~in[141]; 
    assign layer_0[210] = in[346] & in[405]; 
    assign layer_0[211] = in[433] ^ in[660]; 
    assign layer_0[212] = ~(in[292] ^ in[424]); 
    assign layer_0[213] = in[8]; 
    assign layer_0[214] = ~in[481] | (in[75] & in[481]); 
    assign layer_0[215] = ~in[127] | (in[127] & in[654]); 
    assign layer_0[216] = ~(in[326] ^ in[297]); 
    assign layer_0[217] = ~in[628]; 
    assign layer_0[218] = in[248] ^ in[725]; 
    assign layer_0[219] = in[510] & ~in[736]; 
    assign layer_0[220] = ~in[144]; 
    assign layer_0[221] = ~(in[335] & in[438]); 
    assign layer_0[222] = in[507] | in[390]; 
    assign layer_0[223] = in[8] & in[2]; 
    assign layer_0[224] = ~in[585] | (in[262] & in[585]); 
    assign layer_0[225] = in[155] & in[164]; 
    assign layer_0[226] = ~in[237]; 
    assign layer_0[227] = ~(in[609] | in[40]); 
    assign layer_0[228] = in[255] | in[257]; 
    assign layer_0[229] = ~(in[273] | in[441]); 
    assign layer_0[230] = in[675] & in[164]; 
    assign layer_0[231] = in[532] ^ in[339]; 
    assign layer_0[232] = ~(in[485] | in[739]); 
    assign layer_0[233] = in[213] & in[155]; 
    assign layer_0[234] = ~(in[737] | in[347]); 
    assign layer_0[235] = in[761] ^ in[165]; 
    assign layer_0[236] = in[521] & ~in[241]; 
    assign layer_0[237] = in[537] & ~in[744]; 
    assign layer_0[238] = ~in[652] | (in[652] & in[264]); 
    assign layer_0[239] = in[27] ^ in[284]; 
    assign layer_0[240] = ~in[179] | (in[179] & in[435]); 
    assign layer_0[241] = ~in[32] | (in[569] & in[32]); 
    assign layer_0[242] = ~(in[227] ^ in[30]); 
    assign layer_0[243] = in[690] ^ in[697]; 
    assign layer_0[244] = in[321] ^ in[584]; 
    assign layer_0[245] = in[93] & ~in[559]; 
    assign layer_0[246] = in[268] | in[643]; 
    assign layer_0[247] = 1'b1; 
    assign layer_0[248] = in[555] & in[109]; 
    assign layer_0[249] = ~in[255]; 
    assign layer_0[250] = in[608]; 
    assign layer_0[251] = in[665] ^ in[761]; 
    assign layer_0[252] = ~(in[292] ^ in[323]); 
    assign layer_0[253] = in[636] & ~in[520]; 
    assign layer_0[254] = ~(in[375] & in[193]); 
    assign layer_0[255] = ~in[212]; 
    assign layer_0[256] = ~in[316]; 
    assign layer_0[257] = in[370] ^ in[194]; 
    assign layer_0[258] = ~in[109]; 
    assign layer_0[259] = ~(in[251] ^ in[333]); 
    assign layer_0[260] = in[273] ^ in[24]; 
    assign layer_0[261] = in[129]; 
    assign layer_0[262] = ~(in[701] | in[615]); 
    assign layer_0[263] = ~in[227]; 
    assign layer_0[264] = ~(in[453] ^ in[628]); 
    assign layer_0[265] = in[323] ^ in[728]; 
    assign layer_0[266] = ~(in[676] ^ in[599]); 
    assign layer_0[267] = in[328]; 
    assign layer_0[268] = ~in[674]; 
    assign layer_0[269] = in[409] & ~in[357]; 
    assign layer_0[270] = ~in[279]; 
    assign layer_0[271] = ~in[82] | (in[80] & in[82]); 
    assign layer_0[272] = ~(in[633] ^ in[276]); 
    assign layer_0[273] = in[564] | in[500]; 
    assign layer_0[274] = in[616] ^ in[520]; 
    assign layer_0[275] = ~(in[618] ^ in[659]); 
    assign layer_0[276] = ~(in[763] ^ in[754]); 
    assign layer_0[277] = in[503] & ~in[18]; 
    assign layer_0[278] = ~in[249] | (in[541] & in[249]); 
    assign layer_0[279] = ~in[120] | (in[733] & in[120]); 
    assign layer_0[280] = in[131] & ~in[86]; 
    assign layer_0[281] = in[589] | in[669]; 
    assign layer_0[282] = ~in[388] | (in[684] & in[388]); 
    assign layer_0[283] = in[2] ^ in[131]; 
    assign layer_0[284] = ~(in[20] & in[724]); 
    assign layer_0[285] = ~in[158]; 
    assign layer_0[286] = in[469] & ~in[79]; 
    assign layer_0[287] = ~(in[726] & in[173]); 
    assign layer_0[288] = ~(in[533] & in[598]); 
    assign layer_0[289] = in[731] & ~in[141]; 
    assign layer_0[290] = in[265]; 
    assign layer_0[291] = ~(in[146] & in[294]); 
    assign layer_0[292] = in[744] ^ in[712]; 
    assign layer_0[293] = ~in[466]; 
    assign layer_0[294] = ~(in[496] ^ in[285]); 
    assign layer_0[295] = in[451]; 
    assign layer_0[296] = in[379] ^ in[469]; 
    assign layer_0[297] = ~in[474]; 
    assign layer_0[298] = in[35] ^ in[200]; 
    assign layer_0[299] = in[188] | in[289]; 
    assign layer_0[300] = ~in[84]; 
    assign layer_0[301] = ~in[126] | (in[126] & in[219]); 
    assign layer_0[302] = in[243] & ~in[353]; 
    assign layer_0[303] = in[24] & ~in[13]; 
    assign layer_0[304] = in[61] ^ in[482]; 
    assign layer_0[305] = in[646] ^ in[632]; 
    assign layer_0[306] = in[767] & ~in[48]; 
    assign layer_0[307] = ~(in[245] | in[571]); 
    assign layer_0[308] = in[422] ^ in[706]; 
    assign layer_0[309] = ~in[81]; 
    assign layer_0[310] = in[502] ^ in[444]; 
    assign layer_0[311] = in[362] & in[653]; 
    assign layer_0[312] = ~(in[355] ^ in[158]); 
    assign layer_0[313] = in[678] & in[195]; 
    assign layer_0[314] = ~(in[694] ^ in[39]); 
    assign layer_0[315] = ~(in[275] ^ in[664]); 
    assign layer_0[316] = in[52] & ~in[269]; 
    assign layer_0[317] = ~(in[528] | in[324]); 
    assign layer_0[318] = ~(in[251] ^ in[406]); 
    assign layer_0[319] = ~(in[629] & in[237]); 
    assign layer_0[320] = in[13] ^ in[266]; 
    assign layer_0[321] = in[431] & ~in[382]; 
    assign layer_0[322] = ~in[617] | (in[617] & in[668]); 
    assign layer_0[323] = ~(in[131] ^ in[34]); 
    assign layer_0[324] = in[453] ^ in[563]; 
    assign layer_0[325] = ~(in[551] ^ in[760]); 
    assign layer_0[326] = ~in[268] | (in[268] & in[398]); 
    assign layer_0[327] = in[503] & in[295]; 
    assign layer_0[328] = ~in[743]; 
    assign layer_0[329] = ~in[157]; 
    assign layer_0[330] = in[668] ^ in[290]; 
    assign layer_0[331] = ~(in[217] ^ in[319]); 
    assign layer_0[332] = ~(in[307] | in[714]); 
    assign layer_0[333] = in[520] ^ in[522]; 
    assign layer_0[334] = ~(in[36] ^ in[62]); 
    assign layer_0[335] = in[56] ^ in[79]; 
    assign layer_0[336] = in[549] | in[646]; 
    assign layer_0[337] = in[356] ^ in[715]; 
    assign layer_0[338] = in[275] & ~in[447]; 
    assign layer_0[339] = ~in[176]; 
    assign layer_0[340] = in[552] | in[611]; 
    assign layer_0[341] = in[264]; 
    assign layer_0[342] = in[490]; 
    assign layer_0[343] = ~(in[138] & in[520]); 
    assign layer_0[344] = ~(in[582] | in[583]); 
    assign layer_0[345] = ~(in[539] ^ in[506]); 
    assign layer_0[346] = ~in[345] | (in[345] & in[331]); 
    assign layer_0[347] = ~(in[697] ^ in[673]); 
    assign layer_0[348] = in[613] ^ in[745]; 
    assign layer_0[349] = in[173] & ~in[109]; 
    assign layer_0[350] = in[88] & ~in[143]; 
    assign layer_0[351] = in[40] & ~in[607]; 
    assign layer_0[352] = in[550] ^ in[565]; 
    assign layer_0[353] = in[588] & ~in[226]; 
    assign layer_0[354] = ~(in[222] ^ in[492]); 
    assign layer_0[355] = 1'b0; 
    assign layer_0[356] = in[142] & ~in[640]; 
    assign layer_0[357] = ~in[738] | (in[738] & in[113]); 
    assign layer_0[358] = in[177] & ~in[322]; 
    assign layer_0[359] = ~(in[476] & in[92]); 
    assign layer_0[360] = ~(in[700] | in[582]); 
    assign layer_0[361] = in[748] ^ in[555]; 
    assign layer_0[362] = in[28] & in[552]; 
    assign layer_0[363] = in[338] & ~in[370]; 
    assign layer_0[364] = in[613] & ~in[277]; 
    assign layer_0[365] = ~(in[293] & in[504]); 
    assign layer_0[366] = ~(in[745] ^ in[697]); 
    assign layer_0[367] = ~(in[519] & in[242]); 
    assign layer_0[368] = in[375] & in[129]; 
    assign layer_0[369] = ~(in[622] | in[326]); 
    assign layer_0[370] = in[596] & ~in[500]; 
    assign layer_0[371] = in[589] ^ in[332]; 
    assign layer_0[372] = ~(in[637] ^ in[635]); 
    assign layer_0[373] = ~(in[658] | in[682]); 
    assign layer_0[374] = ~(in[760] ^ in[227]); 
    assign layer_0[375] = in[394] & ~in[115]; 
    assign layer_0[376] = in[397] & ~in[22]; 
    assign layer_0[377] = ~in[650] | (in[650] & in[520]); 
    assign layer_0[378] = in[276] & in[709]; 
    assign layer_0[379] = in[411] & ~in[173]; 
    assign layer_0[380] = 1'b0; 
    assign layer_0[381] = ~in[192] | (in[192] & in[371]); 
    assign layer_0[382] = ~in[484]; 
    assign layer_0[383] = ~(in[680] & in[227]); 
    assign layer_0[384] = in[671] & ~in[522]; 
    assign layer_0[385] = in[345] ^ in[413]; 
    assign layer_0[386] = in[96]; 
    assign layer_0[387] = in[334] ^ in[645]; 
    assign layer_0[388] = in[425] & ~in[550]; 
    assign layer_0[389] = in[654] ^ in[28]; 
    assign layer_0[390] = ~(in[632] ^ in[308]); 
    assign layer_0[391] = ~(in[281] ^ in[564]); 
    assign layer_0[392] = ~(in[659] & in[111]); 
    assign layer_0[393] = ~(in[743] ^ in[698]); 
    assign layer_0[394] = ~in[595]; 
    assign layer_0[395] = ~(in[332] & in[651]); 
    assign layer_0[396] = ~(in[282] ^ in[263]); 
    assign layer_0[397] = ~in[574] | (in[574] & in[328]); 
    assign layer_0[398] = in[436]; 
    assign layer_0[399] = ~in[232]; 
    assign layer_0[400] = in[348] & in[603]; 
    assign layer_0[401] = in[621] & ~in[202]; 
    assign layer_0[402] = in[679]; 
    assign layer_0[403] = in[364] & in[44]; 
    assign layer_0[404] = ~(in[483] ^ in[178]); 
    assign layer_0[405] = ~(in[457] ^ in[531]); 
    assign layer_0[406] = in[520] ^ in[622]; 
    assign layer_0[407] = in[652] ^ in[555]; 
    assign layer_0[408] = in[367] ^ in[415]; 
    assign layer_0[409] = in[371] ^ in[153]; 
    assign layer_0[410] = ~(in[297] | in[570]); 
    assign layer_0[411] = in[482] & in[235]; 
    assign layer_0[412] = ~(in[421] | in[467]); 
    assign layer_0[413] = ~(in[583] ^ in[648]); 
    assign layer_0[414] = ~(in[716] ^ in[241]); 
    assign layer_0[415] = ~(in[669] | in[24]); 
    assign layer_0[416] = ~(in[289] | in[258]); 
    assign layer_0[417] = ~in[620] | (in[620] & in[490]); 
    assign layer_0[418] = in[537] ^ in[665]; 
    assign layer_0[419] = ~(in[661] ^ in[664]); 
    assign layer_0[420] = ~(in[587] ^ in[616]); 
    assign layer_0[421] = ~in[299]; 
    assign layer_0[422] = in[726] ^ in[285]; 
    assign layer_0[423] = in[419] & ~in[482]; 
    assign layer_0[424] = in[327]; 
    assign layer_0[425] = ~in[10]; 
    assign layer_0[426] = in[697] ^ in[299]; 
    assign layer_0[427] = ~(in[403] ^ in[386]); 
    assign layer_0[428] = ~(in[667] ^ in[659]); 
    assign layer_0[429] = ~(in[681] & in[372]); 
    assign layer_0[430] = ~(in[690] ^ in[600]); 
    assign layer_0[431] = in[601] ^ in[292]; 
    assign layer_0[432] = in[682] ^ in[649]; 
    assign layer_0[433] = in[92]; 
    assign layer_0[434] = in[758] | in[628]; 
    assign layer_0[435] = 1'b0; 
    assign layer_0[436] = in[647] ^ in[633]; 
    assign layer_0[437] = ~in[395] | (in[395] & in[308]); 
    assign layer_0[438] = in[207] ^ in[78]; 
    assign layer_0[439] = ~(in[658] | in[659]); 
    assign layer_0[440] = ~(in[669] ^ in[70]); 
    assign layer_0[441] = in[197] ^ in[37]; 
    assign layer_0[442] = ~(in[410] & in[646]); 
    assign layer_0[443] = in[646] & ~in[413]; 
    assign layer_0[444] = ~(in[474] ^ in[281]); 
    assign layer_0[445] = ~(in[509] | in[418]); 
    assign layer_0[446] = ~in[487] | (in[688] & in[487]); 
    assign layer_0[447] = in[298] ^ in[613]; 
    assign layer_0[448] = in[588] | in[633]; 
    assign layer_0[449] = ~(in[368] ^ in[206]); 
    assign layer_0[450] = 1'b0; 
    assign layer_0[451] = ~in[486] | (in[754] & in[486]); 
    assign layer_0[452] = ~(in[412] ^ in[446]); 
    assign layer_0[453] = in[63] ^ in[627]; 
    assign layer_0[454] = ~in[579] | (in[579] & in[682]); 
    assign layer_0[455] = ~in[283]; 
    assign layer_0[456] = ~(in[690] ^ in[388]); 
    assign layer_0[457] = in[662] & ~in[641]; 
    assign layer_0[458] = in[567] | in[568]; 
    assign layer_0[459] = in[403] ^ in[193]; 
    assign layer_0[460] = ~(in[553] ^ in[415]); 
    assign layer_0[461] = ~in[445]; 
    assign layer_0[462] = in[325] & ~in[131]; 
    assign layer_0[463] = in[264] & ~in[276]; 
    assign layer_0[464] = ~in[294] | (in[294] & in[694]); 
    assign layer_0[465] = in[507] ^ in[522]; 
    assign layer_0[466] = in[110] | in[262]; 
    assign layer_0[467] = ~in[299]; 
    assign layer_0[468] = in[566]; 
    assign layer_0[469] = ~in[335]; 
    assign layer_0[470] = ~(in[52] | in[610]); 
    assign layer_0[471] = ~(in[730] ^ in[728]); 
    assign layer_0[472] = in[489]; 
    assign layer_0[473] = in[386] | in[109]; 
    assign layer_0[474] = in[179] ^ in[667]; 
    assign layer_0[475] = ~in[662] | (in[36] & in[662]); 
    assign layer_0[476] = ~(in[42] | in[36]); 
    assign layer_0[477] = ~(in[613] ^ in[660]); 
    assign layer_0[478] = in[451] | in[128]; 
    assign layer_0[479] = in[657] ^ in[89]; 
    assign layer_0[480] = ~(in[364] ^ in[702]); 
    assign layer_0[481] = ~(in[103] & in[408]); 
    assign layer_0[482] = in[584] ^ in[205]; 
    assign layer_0[483] = ~(in[686] ^ in[315]); 
    assign layer_0[484] = ~in[505] | (in[227] & in[505]); 
    assign layer_0[485] = ~in[249]; 
    assign layer_0[486] = ~(in[264] | in[725]); 
    assign layer_0[487] = in[89]; 
    assign layer_0[488] = in[695] & in[400]; 
    assign layer_0[489] = in[650] ^ in[70]; 
    assign layer_0[490] = ~(in[365] ^ in[162]); 
    assign layer_0[491] = in[253] | in[668]; 
    assign layer_0[492] = ~in[263] | (in[191] & in[263]); 
    assign layer_0[493] = in[300] & ~in[290]; 
    assign layer_0[494] = ~in[319]; 
    assign layer_0[495] = in[695]; 
    assign layer_0[496] = in[172] & in[375]; 
    assign layer_0[497] = ~(in[297] | in[538]); 
    assign layer_0[498] = in[648]; 
    assign layer_0[499] = in[425] ^ in[565]; 
    assign layer_0[500] = ~(in[714] ^ in[661]); 
    assign layer_0[501] = in[307]; 
    assign layer_0[502] = ~in[332] | (in[656] & in[332]); 
    assign layer_0[503] = in[616] ^ in[631]; 
    assign layer_0[504] = ~(in[73] & in[669]); 
    assign layer_0[505] = in[348] | in[598]; 
    assign layer_0[506] = in[276] ^ in[279]; 
    assign layer_0[507] = in[359] ^ in[261]; 
    assign layer_0[508] = ~in[94] | (in[94] & in[603]); 
    assign layer_0[509] = in[621] & ~in[598]; 
    assign layer_0[510] = ~(in[65] | in[484]); 
    assign layer_0[511] = in[9] & ~in[18]; 
    assign layer_0[512] = ~(in[683] ^ in[617]); 
    assign layer_0[513] = ~in[407]; 
    assign layer_0[514] = in[111] & ~in[746]; 
    assign layer_0[515] = ~in[221]; 
    assign layer_0[516] = ~in[470]; 
    assign layer_0[517] = in[476] ^ in[600]; 
    assign layer_0[518] = in[283] | in[584]; 
    assign layer_0[519] = ~in[683] | (in[227] & in[683]); 
    assign layer_0[520] = in[663] ^ in[226]; 
    assign layer_0[521] = ~(in[261] | in[551]); 
    assign layer_0[522] = ~(in[585] ^ in[566]); 
    assign layer_0[523] = in[195] & in[736]; 
    assign layer_0[524] = ~(in[206] ^ in[381]); 
    assign layer_0[525] = in[171]; 
    assign layer_0[526] = ~(in[19] ^ in[631]); 
    assign layer_0[527] = ~(in[211] | in[625]); 
    assign layer_0[528] = ~(in[576] ^ in[539]); 
    assign layer_0[529] = in[221] & ~in[46]; 
    assign layer_0[530] = ~(in[157] & in[487]); 
    assign layer_0[531] = ~(in[446] | in[46]); 
    assign layer_0[532] = in[95]; 
    assign layer_0[533] = ~in[643]; 
    assign layer_0[534] = in[515] & in[336]; 
    assign layer_0[535] = in[221] & in[53]; 
    assign layer_0[536] = ~in[453] | (in[453] & in[292]); 
    assign layer_0[537] = ~(in[386] | in[340]); 
    assign layer_0[538] = ~(in[74] ^ in[452]); 
    assign layer_0[539] = ~(in[163] ^ in[534]); 
    assign layer_0[540] = ~(in[486] ^ in[183]); 
    assign layer_0[541] = ~in[183] | (in[183] & in[83]); 
    assign layer_0[542] = in[760]; 
    assign layer_0[543] = ~in[397]; 
    assign layer_0[544] = ~in[689]; 
    assign layer_0[545] = in[93] & in[402]; 
    assign layer_0[546] = in[611] ^ in[764]; 
    assign layer_0[547] = ~in[295] | (in[206] & in[295]); 
    assign layer_0[548] = ~in[23] | (in[23] & in[766]); 
    assign layer_0[549] = in[637] & ~in[671]; 
    assign layer_0[550] = in[285] | in[128]; 
    assign layer_0[551] = ~in[282] | (in[282] & in[266]); 
    assign layer_0[552] = ~in[86] | (in[634] & in[86]); 
    assign layer_0[553] = in[697] | in[614]; 
    assign layer_0[554] = ~(in[520] ^ in[693]); 
    assign layer_0[555] = in[493] ^ in[680]; 
    assign layer_0[556] = in[430]; 
    assign layer_0[557] = in[667] ^ in[571]; 
    assign layer_0[558] = in[747]; 
    assign layer_0[559] = in[644] & ~in[613]; 
    assign layer_0[560] = in[710] & ~in[417]; 
    assign layer_0[561] = in[439] | in[500]; 
    assign layer_0[562] = in[324] & ~in[307]; 
    assign layer_0[563] = in[627]; 
    assign layer_0[564] = ~(in[669] | in[518]); 
    assign layer_0[565] = ~(in[54] | in[22]); 
    assign layer_0[566] = ~(in[268] & in[50]); 
    assign layer_0[567] = in[674] ^ in[356]; 
    assign layer_0[568] = ~in[710]; 
    assign layer_0[569] = ~(in[237] ^ in[657]); 
    assign layer_0[570] = ~(in[208] & in[131]); 
    assign layer_0[571] = ~(in[61] | in[539]); 
    assign layer_0[572] = ~in[677]; 
    assign layer_0[573] = ~in[461] | (in[580] & in[461]); 
    assign layer_0[574] = in[688] ^ in[437]; 
    assign layer_0[575] = in[390] | in[328]; 
    assign layer_0[576] = in[418] ^ in[554]; 
    assign layer_0[577] = in[658] | in[208]; 
    assign layer_0[578] = in[139] & ~in[78]; 
    assign layer_0[579] = in[454] & ~in[637]; 
    assign layer_0[580] = in[417] ^ in[609]; 
    assign layer_0[581] = ~in[695] | (in[695] & in[360]); 
    assign layer_0[582] = ~(in[686] ^ in[245]); 
    assign layer_0[583] = in[358] | in[48]; 
    assign layer_0[584] = in[707] | in[612]; 
    assign layer_0[585] = ~(in[229] ^ in[621]); 
    assign layer_0[586] = in[475] ^ in[699]; 
    assign layer_0[587] = in[693] ^ in[83]; 
    assign layer_0[588] = ~(in[427] ^ in[16]); 
    assign layer_0[589] = in[401] & ~in[561]; 
    assign layer_0[590] = ~(in[586] ^ in[585]); 
    assign layer_0[591] = in[548] ^ in[396]; 
    assign layer_0[592] = in[16] | in[524]; 
    assign layer_0[593] = in[141]; 
    assign layer_0[594] = in[631] & ~in[582]; 
    assign layer_0[595] = ~(in[695] | in[658]); 
    assign layer_0[596] = ~in[329]; 
    assign layer_0[597] = ~in[66] | (in[727] & in[66]); 
    assign layer_0[598] = in[147] & ~in[121]; 
    assign layer_0[599] = ~(in[452] & in[61]); 
    assign layer_0[600] = in[534] & ~in[570]; 
    assign layer_0[601] = in[612] & ~in[527]; 
    assign layer_0[602] = in[491] ^ in[568]; 
    assign layer_0[603] = in[94] & in[579]; 
    assign layer_0[604] = ~(in[400] | in[183]); 
    assign layer_0[605] = ~in[311] | (in[311] & in[473]); 
    assign layer_0[606] = in[207] & in[662]; 
    assign layer_0[607] = ~(in[516] | in[50]); 
    assign layer_0[608] = in[387] | in[348]; 
    assign layer_0[609] = ~in[416]; 
    assign layer_0[610] = ~(in[454] ^ in[5]); 
    assign layer_0[611] = ~in[462]; 
    assign layer_0[612] = ~(in[77] ^ in[401]); 
    assign layer_0[613] = in[191] | in[600]; 
    assign layer_0[614] = in[108] | in[568]; 
    assign layer_0[615] = in[371]; 
    assign layer_0[616] = in[715] | in[336]; 
    assign layer_0[617] = in[674]; 
    assign layer_0[618] = ~in[644]; 
    assign layer_0[619] = ~in[206] | (in[206] & in[520]); 
    assign layer_0[620] = in[10] & ~in[666]; 
    assign layer_0[621] = in[648] ^ in[499]; 
    assign layer_0[622] = ~in[24]; 
    assign layer_0[623] = ~in[600] | (in[594] & in[600]); 
    assign layer_0[624] = ~in[23] | (in[23] & in[549]); 
    assign layer_0[625] = 1'b1; 
    assign layer_0[626] = ~in[301]; 
    assign layer_0[627] = ~(in[725] & in[520]); 
    assign layer_0[628] = in[317] & ~in[735]; 
    assign layer_0[629] = ~(in[716] & in[519]); 
    assign layer_0[630] = in[699] | in[519]; 
    assign layer_0[631] = ~in[288]; 
    assign layer_0[632] = 1'b1; 
    assign layer_0[633] = ~in[160]; 
    assign layer_0[634] = in[520] & ~in[488]; 
    assign layer_0[635] = ~(in[662] ^ in[549]); 
    assign layer_0[636] = in[338]; 
    assign layer_0[637] = ~in[51]; 
    assign layer_0[638] = ~(in[277] ^ in[339]); 
    assign layer_0[639] = in[697] & ~in[115]; 
    assign layer_0[640] = ~in[86] | (in[86] & in[321]); 
    assign layer_0[641] = in[367] ^ in[736]; 
    assign layer_0[642] = in[584] ^ in[286]; 
    assign layer_0[643] = ~in[233] | (in[233] & in[100]); 
    assign layer_0[644] = in[436] & ~in[674]; 
    assign layer_0[645] = ~(in[684] & in[518]); 
    assign layer_0[646] = ~(in[319] ^ in[301]); 
    assign layer_0[647] = ~(in[382] ^ in[486]); 
    assign layer_0[648] = in[124] ^ in[482]; 
    assign layer_0[649] = in[678] & in[355]; 
    assign layer_0[650] = ~(in[382] | in[523]); 
    assign layer_0[651] = in[158] & ~in[547]; 
    assign layer_0[652] = in[290]; 
    assign layer_0[653] = ~(in[244] ^ in[110]); 
    assign layer_0[654] = ~in[432]; 
    assign layer_0[655] = in[419]; 
    assign layer_0[656] = ~(in[267] | in[176]); 
    assign layer_0[657] = ~in[144]; 
    assign layer_0[658] = ~in[630]; 
    assign layer_0[659] = in[724] & ~in[32]; 
    assign layer_0[660] = ~in[579] | (in[579] & in[553]); 
    assign layer_0[661] = ~(in[177] | in[539]); 
    assign layer_0[662] = ~in[261]; 
    assign layer_0[663] = ~(in[563] | in[386]); 
    assign layer_0[664] = in[434] & ~in[612]; 
    assign layer_0[665] = in[19] ^ in[398]; 
    assign layer_0[666] = ~in[181] | (in[181] & in[573]); 
    assign layer_0[667] = ~in[678] | (in[678] & in[268]); 
    assign layer_0[668] = in[91] & ~in[27]; 
    assign layer_0[669] = in[76]; 
    assign layer_0[670] = in[181]; 
    assign layer_0[671] = ~(in[484] & in[566]); 
    assign layer_0[672] = in[174] & ~in[375]; 
    assign layer_0[673] = in[215] & ~in[207]; 
    assign layer_0[674] = ~in[568] | (in[568] & in[600]); 
    assign layer_0[675] = in[630] & ~in[444]; 
    assign layer_0[676] = ~(in[413] | in[675]); 
    assign layer_0[677] = ~in[410] | (in[440] & in[410]); 
    assign layer_0[678] = in[614] ^ in[720]; 
    assign layer_0[679] = ~(in[121] & in[288]); 
    assign layer_0[680] = in[185] & ~in[204]; 
    assign layer_0[681] = in[670] ^ in[466]; 
    assign layer_0[682] = in[587] & ~in[761]; 
    assign layer_0[683] = ~(in[484] | in[491]); 
    assign layer_0[684] = in[643] & ~in[328]; 
    assign layer_0[685] = in[667] & in[644]; 
    assign layer_0[686] = in[674] | in[62]; 
    assign layer_0[687] = in[586] & ~in[703]; 
    assign layer_0[688] = in[657] & ~in[653]; 
    assign layer_0[689] = in[3] ^ in[281]; 
    assign layer_0[690] = in[100]; 
    assign layer_0[691] = in[400] & ~in[216]; 
    assign layer_0[692] = ~in[521] | (in[521] & in[555]); 
    assign layer_0[693] = in[556] | in[520]; 
    assign layer_0[694] = ~(in[191] ^ in[684]); 
    assign layer_0[695] = in[686] & ~in[629]; 
    assign layer_0[696] = in[204] ^ in[643]; 
    assign layer_0[697] = ~(in[211] ^ in[569]); 
    assign layer_0[698] = in[571] ^ in[756]; 
    assign layer_0[699] = ~(in[645] ^ in[583]); 
    assign layer_0[700] = in[264] ^ in[282]; 
    assign layer_0[701] = in[727] | in[701]; 
    assign layer_0[702] = ~(in[535] ^ in[508]); 
    assign layer_0[703] = in[315] & ~in[207]; 
    assign layer_0[704] = ~(in[600] ^ in[554]); 
    assign layer_0[705] = ~in[504] | (in[504] & in[140]); 
    assign layer_0[706] = in[298] & ~in[761]; 
    assign layer_0[707] = ~in[282] | (in[5] & in[282]); 
    assign layer_0[708] = in[604] ^ in[562]; 
    assign layer_0[709] = in[747] & ~in[744]; 
    assign layer_0[710] = ~(in[263] | in[681]); 
    assign layer_0[711] = in[156] ^ in[637]; 
    assign layer_0[712] = ~in[533]; 
    assign layer_0[713] = ~in[379] | (in[490] & in[379]); 
    assign layer_0[714] = ~in[302] | (in[302] & in[417]); 
    assign layer_0[715] = in[741] & ~in[512]; 
    assign layer_0[716] = in[397] & in[416]; 
    assign layer_0[717] = in[743]; 
    assign layer_0[718] = in[250] & ~in[731]; 
    assign layer_0[719] = in[353] | in[490]; 
    assign layer_0[720] = in[666] | in[3]; 
    assign layer_0[721] = in[311] ^ in[489]; 
    assign layer_0[722] = in[741] & ~in[14]; 
    assign layer_0[723] = ~(in[126] | in[469]); 
    assign layer_0[724] = in[226] ^ in[97]; 
    assign layer_0[725] = in[388] ^ in[688]; 
    assign layer_0[726] = ~(in[743] & in[151]); 
    assign layer_0[727] = in[655] ^ in[710]; 
    assign layer_0[728] = ~in[145]; 
    assign layer_0[729] = ~in[328] | (in[296] & in[328]); 
    assign layer_0[730] = ~in[173]; 
    assign layer_0[731] = ~in[539]; 
    assign layer_0[732] = ~(in[13] ^ in[423]); 
    assign layer_0[733] = ~in[119] | (in[119] & in[715]); 
    assign layer_0[734] = ~in[350] | (in[210] & in[350]); 
    assign layer_0[735] = in[414] & ~in[422]; 
    assign layer_0[736] = in[645] & in[435]; 
    assign layer_0[737] = in[395]; 
    assign layer_0[738] = ~(in[455] ^ in[764]); 
    assign layer_0[739] = ~(in[298] | in[44]); 
    assign layer_0[740] = ~(in[388] ^ in[710]); 
    assign layer_0[741] = in[744]; 
    assign layer_0[742] = in[603] & ~in[232]; 
    assign layer_0[743] = ~(in[699] | in[388]); 
    assign layer_0[744] = in[67] ^ in[209]; 
    assign layer_0[745] = ~in[713]; 
    assign layer_0[746] = in[149] & ~in[324]; 
    assign layer_0[747] = in[571]; 
    assign layer_0[748] = in[520] & in[518]; 
    assign layer_0[749] = in[697] ^ in[492]; 
    assign layer_0[750] = in[618] ^ in[318]; 
    assign layer_0[751] = ~(in[569] ^ in[552]); 
    assign layer_0[752] = ~(in[509] & in[534]); 
    assign layer_0[753] = in[180] ^ in[451]; 
    assign layer_0[754] = ~(in[697] & in[131]); 
    assign layer_0[755] = in[587] ^ in[40]; 
    assign layer_0[756] = in[55] & ~in[508]; 
    assign layer_0[757] = in[250] | in[715]; 
    assign layer_0[758] = in[250]; 
    assign layer_0[759] = in[649] & ~in[386]; 
    assign layer_0[760] = in[342] | in[681]; 
    assign layer_0[761] = ~in[43] | (in[565] & in[43]); 
    assign layer_0[762] = in[104] & in[292]; 
    assign layer_0[763] = in[612] | in[649]; 
    assign layer_0[764] = in[746]; 
    assign layer_0[765] = ~(in[334] ^ in[659]); 
    assign layer_0[766] = in[707] ^ in[307]; 
    assign layer_0[767] = in[212]; 
    assign layer_0[768] = ~in[691]; 
    assign layer_0[769] = in[233] & ~in[545]; 
    assign layer_0[770] = ~in[327] | (in[327] & in[600]); 
    assign layer_0[771] = in[18] ^ in[488]; 
    assign layer_0[772] = in[172] & in[602]; 
    assign layer_0[773] = ~(in[536] ^ in[28]); 
    assign layer_0[774] = ~in[354] | (in[354] & in[271]); 
    assign layer_0[775] = ~(in[61] ^ in[115]); 
    assign layer_0[776] = ~(in[584] & in[25]); 
    assign layer_0[777] = in[381]; 
    assign layer_0[778] = in[647] & ~in[177]; 
    assign layer_0[779] = in[431] | in[38]; 
    assign layer_0[780] = ~in[682]; 
    assign layer_0[781] = in[204]; 
    assign layer_0[782] = ~in[109] | (in[54] & in[109]); 
    assign layer_0[783] = in[252]; 
    assign layer_0[784] = in[606] ^ in[639]; 
    assign layer_0[785] = ~(in[78] & in[94]); 
    assign layer_0[786] = in[585] ^ in[491]; 
    assign layer_0[787] = ~(in[318] | in[277]); 
    assign layer_0[788] = in[622]; 
    assign layer_0[789] = in[553]; 
    assign layer_0[790] = in[360]; 
    assign layer_0[791] = in[619]; 
    assign layer_0[792] = in[371]; 
    assign layer_0[793] = in[22] & in[236]; 
    assign layer_0[794] = ~in[549]; 
    assign layer_0[795] = in[12]; 
    assign layer_0[796] = ~(in[588] | in[553]); 
    assign layer_0[797] = ~(in[128] & in[348]); 
    assign layer_0[798] = ~in[37]; 
    assign layer_0[799] = ~in[713] | (in[713] & in[708]); 
    assign layer_0[800] = ~in[318] | (in[646] & in[318]); 
    assign layer_0[801] = ~(in[555] | in[528]); 
    assign layer_0[802] = in[291] ^ in[253]; 
    assign layer_0[803] = ~(in[190] | in[463]); 
    assign layer_0[804] = ~(in[631] | in[539]); 
    assign layer_0[805] = ~in[19]; 
    assign layer_0[806] = in[419] & in[686]; 
    assign layer_0[807] = in[243] | in[253]; 
    assign layer_0[808] = ~in[669] | (in[85] & in[669]); 
    assign layer_0[809] = ~(in[1] | in[378]); 
    assign layer_0[810] = ~(in[617] ^ in[252]); 
    assign layer_0[811] = in[603] & ~in[470]; 
    assign layer_0[812] = in[247]; 
    assign layer_0[813] = in[93] & in[418]; 
    assign layer_0[814] = ~(in[612] ^ in[603]); 
    assign layer_0[815] = ~(in[712] ^ in[714]); 
    assign layer_0[816] = ~(in[537] ^ in[249]); 
    assign layer_0[817] = in[424] & ~in[661]; 
    assign layer_0[818] = in[518] & in[360]; 
    assign layer_0[819] = in[369] ^ in[606]; 
    assign layer_0[820] = in[61] & ~in[584]; 
    assign layer_0[821] = ~in[748] | (in[607] & in[748]); 
    assign layer_0[822] = ~in[396] | (in[396] & in[512]); 
    assign layer_0[823] = in[715] ^ in[439]; 
    assign layer_0[824] = in[160] & ~in[43]; 
    assign layer_0[825] = in[34]; 
    assign layer_0[826] = in[639] & in[639]; 
    assign layer_0[827] = ~in[448] | (in[448] & in[750]); 
    assign layer_0[828] = ~(in[638] ^ in[424]); 
    assign layer_0[829] = in[319] | in[339]; 
    assign layer_0[830] = in[178] | in[475]; 
    assign layer_0[831] = in[584] & ~in[336]; 
    assign layer_0[832] = in[516]; 
    assign layer_0[833] = in[140]; 
    assign layer_0[834] = in[345]; 
    assign layer_0[835] = in[229] & in[557]; 
    assign layer_0[836] = ~in[345]; 
    assign layer_0[837] = ~in[363] | (in[363] & in[66]); 
    assign layer_0[838] = ~(in[606] ^ in[154]); 
    assign layer_0[839] = ~(in[280] ^ in[256]); 
    assign layer_0[840] = ~(in[516] | in[174]); 
    assign layer_0[841] = ~(in[215] ^ in[626]); 
    assign layer_0[842] = ~(in[532] | in[741]); 
    assign layer_0[843] = in[693] | in[568]; 
    assign layer_0[844] = in[126] ^ in[371]; 
    assign layer_0[845] = ~(in[531] ^ in[702]); 
    assign layer_0[846] = ~in[476] | (in[476] & in[631]); 
    assign layer_0[847] = in[141] | in[667]; 
    assign layer_0[848] = in[471]; 
    assign layer_0[849] = ~(in[663] ^ in[416]); 
    assign layer_0[850] = ~in[490]; 
    assign layer_0[851] = ~in[569] | (in[629] & in[569]); 
    assign layer_0[852] = in[651] & ~in[580]; 
    assign layer_0[853] = in[722] ^ in[573]; 
    assign layer_0[854] = in[518] ^ in[650]; 
    assign layer_0[855] = ~in[445] | (in[543] & in[445]); 
    assign layer_0[856] = ~in[282]; 
    assign layer_0[857] = ~in[133]; 
    assign layer_0[858] = ~(in[298] & in[52]); 
    assign layer_0[859] = in[486] ^ in[114]; 
    assign layer_0[860] = ~in[399] | (in[399] & in[10]); 
    assign layer_0[861] = ~(in[651] & in[697]); 
    assign layer_0[862] = in[47] & ~in[36]; 
    assign layer_0[863] = ~(in[342] ^ in[630]); 
    assign layer_0[864] = ~(in[29] ^ in[238]); 
    assign layer_0[865] = in[579]; 
    assign layer_0[866] = in[130] & ~in[551]; 
    assign layer_0[867] = in[376]; 
    assign layer_0[868] = ~in[79] | (in[79] & in[17]); 
    assign layer_0[869] = in[11]; 
    assign layer_0[870] = ~in[423] | (in[387] & in[423]); 
    assign layer_0[871] = ~(in[708] ^ in[557]); 
    assign layer_0[872] = ~(in[421] ^ in[124]); 
    assign layer_0[873] = ~(in[5] ^ in[657]); 
    assign layer_0[874] = in[12] ^ in[743]; 
    assign layer_0[875] = in[293] ^ in[402]; 
    assign layer_0[876] = in[475] & ~in[568]; 
    assign layer_0[877] = ~in[315]; 
    assign layer_0[878] = in[414] | in[710]; 
    assign layer_0[879] = ~in[370]; 
    assign layer_0[880] = ~(in[554] | in[725]); 
    assign layer_0[881] = in[650] & ~in[596]; 
    assign layer_0[882] = ~in[598] | (in[364] & in[598]); 
    assign layer_0[883] = in[561] ^ in[408]; 
    assign layer_0[884] = in[387] & ~in[609]; 
    assign layer_0[885] = in[444] | in[240]; 
    assign layer_0[886] = in[712] & ~in[267]; 
    assign layer_0[887] = ~in[678] | (in[627] & in[678]); 
    assign layer_0[888] = ~in[618] | (in[618] & in[330]); 
    assign layer_0[889] = ~(in[474] ^ in[495]); 
    assign layer_0[890] = ~(in[530] | in[686]); 
    assign layer_0[891] = ~in[98] | (in[5] & in[98]); 
    assign layer_0[892] = ~(in[367] ^ in[533]); 
    assign layer_0[893] = in[263] ^ in[18]; 
    assign layer_0[894] = ~(in[94] | in[156]); 
    assign layer_0[895] = ~in[48]; 
    assign layer_0[896] = in[327] | in[527]; 
    assign layer_0[897] = ~(in[504] & in[152]); 
    assign layer_0[898] = in[253] & ~in[329]; 
    assign layer_0[899] = in[521] | in[396]; 
    assign layer_0[900] = in[262]; 
    assign layer_0[901] = ~(in[626] ^ in[227]); 
    assign layer_0[902] = ~(in[420] | in[66]); 
    assign layer_0[903] = in[477] | in[27]; 
    assign layer_0[904] = ~in[572] | (in[237] & in[572]); 
    assign layer_0[905] = ~in[605] | (in[605] & in[627]); 
    assign layer_0[906] = in[601] & in[136]; 
    assign layer_0[907] = in[418] & ~in[456]; 
    assign layer_0[908] = in[66] | in[596]; 
    assign layer_0[909] = ~in[83] | (in[83] & in[518]); 
    assign layer_0[910] = in[117] | in[609]; 
    assign layer_0[911] = ~(in[325] ^ in[552]); 
    assign layer_0[912] = ~in[13]; 
    assign layer_0[913] = ~(in[3] & in[370]); 
    assign layer_0[914] = ~(in[666] ^ in[379]); 
    assign layer_0[915] = in[305] | in[525]; 
    assign layer_0[916] = in[207]; 
    assign layer_0[917] = ~in[752]; 
    assign layer_0[918] = in[400]; 
    assign layer_0[919] = ~(in[552] ^ in[553]); 
    assign layer_0[920] = ~in[268] | (in[268] & in[623]); 
    assign layer_0[921] = in[26]; 
    assign layer_0[922] = ~in[280]; 
    assign layer_0[923] = in[279]; 
    assign layer_0[924] = in[633]; 
    assign layer_0[925] = in[475] ^ in[586]; 
    assign layer_0[926] = in[697] ^ in[227]; 
    assign layer_0[927] = ~in[391]; 
    assign layer_0[928] = in[550] | in[549]; 
    assign layer_0[929] = in[585]; 
    assign layer_0[930] = in[699] ^ in[570]; 
    assign layer_0[931] = ~in[188] | (in[526] & in[188]); 
    assign layer_0[932] = ~in[622] | (in[26] & in[622]); 
    assign layer_0[933] = in[467] & ~in[299]; 
    assign layer_0[934] = ~(in[693] ^ in[554]); 
    assign layer_0[935] = in[289] ^ in[665]; 
    assign layer_0[936] = ~(in[647] ^ in[649]); 
    assign layer_0[937] = ~(in[233] | in[97]); 
    assign layer_0[938] = ~in[680]; 
    assign layer_0[939] = ~(in[330] ^ in[492]); 
    assign layer_0[940] = ~in[725] | (in[725] & in[472]); 
    assign layer_0[941] = ~(in[415] | in[483]); 
    assign layer_0[942] = ~in[420] | (in[420] & in[516]); 
    assign layer_0[943] = in[378] ^ in[405]; 
    assign layer_0[944] = in[486] ^ in[518]; 
    assign layer_0[945] = in[312] | in[258]; 
    assign layer_0[946] = in[571] ^ in[192]; 
    assign layer_0[947] = ~(in[466] ^ in[332]); 
    assign layer_0[948] = in[718] ^ in[318]; 
    assign layer_0[949] = ~(in[685] | in[284]); 
    assign layer_0[950] = in[399] & ~in[214]; 
    assign layer_0[951] = in[630]; 
    assign layer_0[952] = ~(in[123] & in[647]); 
    assign layer_0[953] = in[531] & ~in[373]; 
    assign layer_0[954] = in[334] & in[111]; 
    assign layer_0[955] = ~in[63] | (in[63] & in[463]); 
    assign layer_0[956] = ~(in[219] ^ in[697]); 
    assign layer_0[957] = in[439]; 
    assign layer_0[958] = in[101] & in[587]; 
    assign layer_0[959] = ~in[651]; 
    assign layer_0[960] = ~(in[665] ^ in[12]); 
    assign layer_0[961] = in[247]; 
    assign layer_0[962] = in[635] ^ in[174]; 
    assign layer_0[963] = ~(in[418] ^ in[693]); 
    assign layer_0[964] = ~(in[338] ^ in[692]); 
    assign layer_0[965] = in[262] | in[651]; 
    assign layer_0[966] = ~(in[323] | in[179]); 
    assign layer_0[967] = ~(in[460] ^ in[696]); 
    assign layer_0[968] = ~(in[210] ^ in[657]); 
    assign layer_0[969] = ~(in[354] ^ in[680]); 
    assign layer_0[970] = ~(in[600] | in[614]); 
    assign layer_0[971] = ~(in[387] | in[683]); 
    assign layer_0[972] = in[40]; 
    assign layer_0[973] = in[8] & in[359]; 
    assign layer_0[974] = in[709] ^ in[206]; 
    assign layer_0[975] = in[694]; 
    assign layer_0[976] = ~in[18]; 
    assign layer_0[977] = ~in[442] | (in[442] & in[482]); 
    assign layer_0[978] = in[759] ^ in[262]; 
    assign layer_0[979] = in[72]; 
    assign layer_0[980] = in[251] | in[647]; 
    assign layer_0[981] = ~in[554]; 
    assign layer_0[982] = ~in[341]; 
    assign layer_0[983] = in[424] ^ in[81]; 
    assign layer_0[984] = ~in[624]; 
    assign layer_0[985] = in[433]; 
    assign layer_0[986] = ~(in[646] ^ in[598]); 
    assign layer_0[987] = ~(in[503] ^ in[3]); 
    assign layer_0[988] = in[277] & ~in[398]; 
    assign layer_0[989] = ~(in[650] ^ in[621]); 
    assign layer_0[990] = in[741] & in[253]; 
    assign layer_0[991] = 1'b0; 
    assign layer_0[992] = ~(in[12] ^ in[261]); 
    assign layer_0[993] = in[695] & ~in[450]; 
    assign layer_0[994] = in[238] | in[535]; 
    assign layer_0[995] = in[205] ^ in[655]; 
    assign layer_0[996] = ~(in[243] ^ in[502]); 
    assign layer_0[997] = in[103] & in[313]; 
    assign layer_0[998] = in[195]; 
    assign layer_0[999] = in[381] & ~in[637]; 
    assign layer_0[1000] = ~(in[731] ^ in[682]); 
    assign layer_0[1001] = ~in[485]; 
    assign layer_0[1002] = in[412] & ~in[596]; 
    assign layer_0[1003] = ~in[230]; 
    assign layer_0[1004] = ~(in[403] ^ in[613]); 
    assign layer_0[1005] = in[714] & in[580]; 
    assign layer_0[1006] = ~(in[239] | in[584]); 
    assign layer_0[1007] = in[765]; 
    assign layer_0[1008] = ~(in[331] ^ in[95]); 
    assign layer_0[1009] = ~(in[324] & in[468]); 
    assign layer_0[1010] = in[25] ^ in[615]; 
    assign layer_0[1011] = ~in[710] | (in[742] & in[710]); 
    assign layer_0[1012] = ~(in[673] ^ in[201]); 
    assign layer_0[1013] = ~(in[599] ^ in[354]); 
    assign layer_0[1014] = in[623] ^ in[341]; 
    assign layer_0[1015] = in[600] ^ in[420]; 
    assign layer_0[1016] = in[304] ^ in[251]; 
    assign layer_0[1017] = ~(in[576] ^ in[151]); 
    assign layer_0[1018] = in[564] ^ in[14]; 
    assign layer_0[1019] = ~(in[10] & in[194]); 
    assign layer_0[1020] = ~(in[628] ^ in[465]); 
    assign layer_0[1021] = ~in[236] | (in[236] & in[361]); 
    assign layer_0[1022] = ~(in[367] & in[235]); 
    assign layer_0[1023] = in[563] & ~in[609]; 
    assign layer_0[1024] = ~(in[345] ^ in[210]); 
    assign layer_0[1025] = in[292] ^ in[487]; 
    assign layer_0[1026] = ~(in[421] ^ in[734]); 
    assign layer_0[1027] = in[469] & in[310]; 
    assign layer_0[1028] = ~(in[501] & in[729]); 
    assign layer_0[1029] = ~in[472] | (in[597] & in[472]); 
    assign layer_0[1030] = in[628]; 
    assign layer_0[1031] = in[34]; 
    assign layer_0[1032] = in[686] | in[697]; 
    assign layer_0[1033] = 1'b1; 
    assign layer_0[1034] = in[75] ^ in[554]; 
    assign layer_0[1035] = ~(in[719] | in[571]); 
    assign layer_0[1036] = ~(in[635] | in[235]); 
    assign layer_0[1037] = in[49] ^ in[366]; 
    assign layer_0[1038] = in[758] ^ in[428]; 
    assign layer_0[1039] = ~in[428] | (in[428] & in[263]); 
    assign layer_0[1040] = ~in[74]; 
    assign layer_0[1041] = ~in[5]; 
    assign layer_0[1042] = in[672] ^ in[379]; 
    assign layer_0[1043] = ~in[82]; 
    assign layer_0[1044] = ~(in[81] ^ in[194]); 
    assign layer_0[1045] = ~in[553] | (in[741] & in[553]); 
    assign layer_0[1046] = in[251]; 
    assign layer_0[1047] = ~(in[388] ^ in[45]); 
    assign layer_0[1048] = in[605] ^ in[277]; 
    assign layer_0[1049] = ~(in[641] ^ in[628]); 
    assign layer_0[1050] = ~(in[445] & in[110]); 
    assign layer_0[1051] = in[616] ^ in[690]; 
    assign layer_0[1052] = in[142] ^ in[335]; 
    assign layer_0[1053] = ~(in[711] & in[239]); 
    assign layer_0[1054] = in[238] ^ in[483]; 
    assign layer_0[1055] = in[358]; 
    assign layer_0[1056] = ~(in[678] ^ in[586]); 
    assign layer_0[1057] = ~(in[45] ^ in[443]); 
    assign layer_0[1058] = ~(in[76] | in[521]); 
    assign layer_0[1059] = ~in[324]; 
    assign layer_0[1060] = in[544] & ~in[26]; 
    assign layer_0[1061] = in[645] & ~in[210]; 
    assign layer_0[1062] = ~(in[354] ^ in[263]); 
    assign layer_0[1063] = in[217] & ~in[367]; 
    assign layer_0[1064] = 1'b1; 
    assign layer_0[1065] = ~in[253]; 
    assign layer_0[1066] = ~(in[304] | in[743]); 
    assign layer_0[1067] = in[39] & ~in[611]; 
    assign layer_0[1068] = ~in[424]; 
    assign layer_0[1069] = in[300] | in[503]; 
    assign layer_0[1070] = in[280] & in[403]; 
    assign layer_0[1071] = ~in[72] | (in[279] & in[72]); 
    assign layer_0[1072] = ~(in[486] ^ in[659]); 
    assign layer_0[1073] = in[506]; 
    assign layer_0[1074] = ~in[672] | (in[196] & in[672]); 
    assign layer_0[1075] = in[582] ^ in[568]; 
    assign layer_0[1076] = in[371] ^ in[244]; 
    assign layer_0[1077] = in[62] ^ in[101]; 
    assign layer_0[1078] = ~(in[355] ^ in[359]); 
    assign layer_0[1079] = ~in[165] | (in[644] & in[165]); 
    assign layer_0[1080] = ~(in[32] ^ in[27]); 
    assign layer_0[1081] = ~in[573] | (in[455] & in[573]); 
    assign layer_0[1082] = ~in[189] | (in[176] & in[189]); 
    assign layer_0[1083] = ~in[438] | (in[438] & in[544]); 
    assign layer_0[1084] = ~in[360]; 
    assign layer_0[1085] = ~(in[410] ^ in[134]); 
    assign layer_0[1086] = in[682] ^ in[664]; 
    assign layer_0[1087] = in[260] ^ in[93]; 
    assign layer_0[1088] = ~(in[317] | in[32]); 
    assign layer_0[1089] = in[568]; 
    assign layer_0[1090] = ~(in[350] & in[161]); 
    assign layer_0[1091] = ~(in[362] ^ in[616]); 
    assign layer_0[1092] = in[717] & ~in[44]; 
    assign layer_0[1093] = ~in[491]; 
    assign layer_0[1094] = 1'b0; 
    assign layer_0[1095] = in[555] ^ in[664]; 
    assign layer_0[1096] = in[491] | in[506]; 
    assign layer_0[1097] = ~(in[222] ^ in[201]); 
    assign layer_0[1098] = ~in[551] | (in[97] & in[551]); 
    assign layer_0[1099] = in[623] & in[600]; 
    assign layer_0[1100] = ~(in[684] ^ in[77]); 
    assign layer_0[1101] = ~in[130]; 
    assign layer_0[1102] = ~in[378] | (in[378] & in[751]); 
    assign layer_0[1103] = in[234] ^ in[702]; 
    assign layer_0[1104] = ~in[126] | (in[644] & in[126]); 
    assign layer_0[1105] = in[43] | in[614]; 
    assign layer_0[1106] = in[569] & ~in[28]; 
    assign layer_0[1107] = ~in[694] | (in[668] & in[694]); 
    assign layer_0[1108] = in[343] ^ in[601]; 
    assign layer_0[1109] = in[24] ^ in[477]; 
    assign layer_0[1110] = ~(in[432] ^ in[217]); 
    assign layer_0[1111] = ~(in[472] ^ in[674]); 
    assign layer_0[1112] = ~(in[310] & in[731]); 
    assign layer_0[1113] = ~in[329]; 
    assign layer_0[1114] = in[351] ^ in[362]; 
    assign layer_0[1115] = in[111]; 
    assign layer_0[1116] = in[672] ^ in[341]; 
    assign layer_0[1117] = ~(in[533] ^ in[549]); 
    assign layer_0[1118] = in[280] ^ in[189]; 
    assign layer_0[1119] = in[161] & in[229]; 
    assign layer_0[1120] = in[339] ^ in[403]; 
    assign layer_0[1121] = ~in[533]; 
    assign layer_0[1122] = in[507] | in[66]; 
    assign layer_0[1123] = ~(in[277] ^ in[569]); 
    assign layer_0[1124] = ~(in[667] ^ in[261]); 
    assign layer_0[1125] = in[522] ^ in[548]; 
    assign layer_0[1126] = in[116] ^ in[669]; 
    assign layer_0[1127] = ~in[296] | (in[296] & in[266]); 
    assign layer_0[1128] = in[521] ^ in[447]; 
    assign layer_0[1129] = in[684] & in[636]; 
    assign layer_0[1130] = ~in[697] | (in[338] & in[697]); 
    assign layer_0[1131] = ~in[379] | (in[679] & in[379]); 
    assign layer_0[1132] = in[662] ^ in[664]; 
    assign layer_0[1133] = ~(in[4] ^ in[61]); 
    assign layer_0[1134] = in[732] ^ in[326]; 
    assign layer_0[1135] = ~(in[137] ^ in[507]); 
    assign layer_0[1136] = ~in[521] | (in[90] & in[521]); 
    assign layer_0[1137] = in[716] | in[45]; 
    assign layer_0[1138] = ~in[461] | (in[210] & in[461]); 
    assign layer_0[1139] = ~in[680]; 
    assign layer_0[1140] = in[278] & ~in[499]; 
    assign layer_0[1141] = ~(in[759] & in[435]); 
    assign layer_0[1142] = in[473] ^ in[338]; 
    assign layer_0[1143] = ~in[682] | (in[682] & in[355]); 
    assign layer_0[1144] = in[733] & ~in[384]; 
    assign layer_0[1145] = ~(in[262] ^ in[263]); 
    assign layer_0[1146] = ~(in[325] & in[243]); 
    assign layer_0[1147] = ~(in[324] ^ in[36]); 
    assign layer_0[1148] = ~(in[61] | in[569]); 
    assign layer_0[1149] = in[730]; 
    assign layer_0[1150] = in[426] & ~in[728]; 
    assign layer_0[1151] = in[361] & in[248]; 
    assign layer_0[1152] = in[615] & ~in[650]; 
    assign layer_0[1153] = ~(in[679] ^ in[643]); 
    assign layer_0[1154] = ~in[456] | (in[132] & in[456]); 
    assign layer_0[1155] = ~in[129]; 
    assign layer_0[1156] = in[631] ^ in[603]; 
    assign layer_0[1157] = in[411] & ~in[741]; 
    assign layer_0[1158] = ~(in[495] ^ in[521]); 
    assign layer_0[1159] = ~(in[739] | in[450]); 
    assign layer_0[1160] = in[602] ^ in[538]; 
    assign layer_0[1161] = ~in[635] | (in[635] & in[440]); 
    assign layer_0[1162] = in[585] ^ in[584]; 
    assign layer_0[1163] = ~(in[362] ^ in[751]); 
    assign layer_0[1164] = in[451]; 
    assign layer_0[1165] = ~(in[205] ^ in[355]); 
    assign layer_0[1166] = ~in[681] | (in[267] & in[681]); 
    assign layer_0[1167] = ~in[501]; 
    assign layer_0[1168] = in[332] & ~in[596]; 
    assign layer_0[1169] = in[308] & in[243]; 
    assign layer_0[1170] = ~(in[760] ^ in[212]); 
    assign layer_0[1171] = in[500] ^ in[327]; 
    assign layer_0[1172] = ~in[128] | (in[128] & in[715]); 
    assign layer_0[1173] = in[680] | in[254]; 
    assign layer_0[1174] = in[391] & ~in[262]; 
    assign layer_0[1175] = in[340] | in[583]; 
    assign layer_0[1176] = in[405] & ~in[466]; 
    assign layer_0[1177] = in[709] ^ in[200]; 
    assign layer_0[1178] = ~(in[676] ^ in[500]); 
    assign layer_0[1179] = ~in[565] | (in[713] & in[565]); 
    assign layer_0[1180] = ~in[474] | (in[236] & in[474]); 
    assign layer_0[1181] = in[551]; 
    assign layer_0[1182] = in[340] ^ in[759]; 
    assign layer_0[1183] = ~(in[12] | in[45]); 
    assign layer_0[1184] = ~in[676] | (in[391] & in[676]); 
    assign layer_0[1185] = in[634] ^ in[618]; 
    assign layer_0[1186] = ~(in[746] | in[385]); 
    assign layer_0[1187] = ~in[421]; 
    assign layer_0[1188] = in[103] & in[407]; 
    assign layer_0[1189] = in[629]; 
    assign layer_0[1190] = in[334] ^ in[421]; 
    assign layer_0[1191] = ~(in[740] ^ in[403]); 
    assign layer_0[1192] = ~(in[170] ^ in[8]); 
    assign layer_0[1193] = in[231] & in[69]; 
    assign layer_0[1194] = in[508] & ~in[305]; 
    assign layer_0[1195] = ~(in[435] | in[760]); 
    assign layer_0[1196] = ~in[450]; 
    assign layer_0[1197] = in[632] & ~in[556]; 
    assign layer_0[1198] = ~(in[502] & in[147]); 
    assign layer_0[1199] = ~(in[305] & in[113]); 
    assign layer_0[1200] = in[619] ^ in[744]; 
    assign layer_0[1201] = ~in[445] | (in[445] & in[486]); 
    assign layer_0[1202] = in[317] & ~in[620]; 
    assign layer_0[1203] = ~in[436] | (in[436] & in[589]); 
    assign layer_0[1204] = in[227] ^ in[622]; 
    assign layer_0[1205] = in[603]; 
    assign layer_0[1206] = in[70] ^ in[588]; 
    assign layer_0[1207] = in[522] ^ in[378]; 
    assign layer_0[1208] = ~in[411] | (in[449] & in[411]); 
    assign layer_0[1209] = ~(in[355] ^ in[731]); 
    assign layer_0[1210] = ~(in[563] & in[656]); 
    assign layer_0[1211] = ~in[137] | (in[22] & in[137]); 
    assign layer_0[1212] = ~(in[555] | in[211]); 
    assign layer_0[1213] = in[630] & ~in[207]; 
    assign layer_0[1214] = in[55] | in[721]; 
    assign layer_0[1215] = in[345] ^ in[755]; 
    assign layer_0[1216] = ~(in[206] ^ in[572]); 
    assign layer_0[1217] = 1'b0; 
    assign layer_0[1218] = ~(in[21] & in[372]); 
    assign layer_0[1219] = ~in[293]; 
    assign layer_0[1220] = in[548] ^ in[307]; 
    assign layer_0[1221] = ~in[182] | (in[127] & in[182]); 
    assign layer_0[1222] = ~in[473] | (in[195] & in[473]); 
    assign layer_0[1223] = in[76] ^ in[275]; 
    assign layer_0[1224] = in[537] ^ in[267]; 
    assign layer_0[1225] = in[175] | in[663]; 
    assign layer_0[1226] = ~in[222]; 
    assign layer_0[1227] = ~in[352] | (in[302] & in[352]); 
    assign layer_0[1228] = in[444] & in[361]; 
    assign layer_0[1229] = ~in[443] | (in[443] & in[288]); 
    assign layer_0[1230] = in[569] & ~in[492]; 
    assign layer_0[1231] = ~(in[416] ^ in[536]); 
    assign layer_0[1232] = ~(in[252] | in[538]); 
    assign layer_0[1233] = in[397] | in[537]; 
    assign layer_0[1234] = ~(in[388] ^ in[746]); 
    assign layer_0[1235] = ~in[677] | (in[677] & in[270]); 
    assign layer_0[1236] = in[341] & ~in[128]; 
    assign layer_0[1237] = ~(in[458] & in[457]); 
    assign layer_0[1238] = ~(in[632] | in[291]); 
    assign layer_0[1239] = 1'b0; 
    assign layer_0[1240] = in[227] & ~in[420]; 
    assign layer_0[1241] = in[315] & ~in[282]; 
    assign layer_0[1242] = ~in[509]; 
    assign layer_0[1243] = ~(in[473] | in[613]); 
    assign layer_0[1244] = ~(in[445] & in[299]); 
    assign layer_0[1245] = in[324] & ~in[592]; 
    assign layer_0[1246] = ~(in[348] | in[673]); 
    assign layer_0[1247] = ~in[507] | (in[476] & in[507]); 
    assign layer_0[1248] = in[538] ^ in[713]; 
    assign layer_0[1249] = in[425] | in[475]; 
    assign layer_0[1250] = ~(in[94] ^ in[325]); 
    assign layer_0[1251] = in[456] & ~in[650]; 
    assign layer_0[1252] = ~in[276] | (in[276] & in[397]); 
    assign layer_0[1253] = in[662] & ~in[628]; 
    assign layer_0[1254] = in[708] | in[307]; 
    assign layer_0[1255] = in[631] & ~in[668]; 
    assign layer_0[1256] = ~(in[733] | in[733]); 
    assign layer_0[1257] = in[53] | in[575]; 
    assign layer_0[1258] = 1'b1; 
    assign layer_0[1259] = in[472]; 
    assign layer_0[1260] = in[98]; 
    assign layer_0[1261] = ~(in[682] | in[475]); 
    assign layer_0[1262] = in[456] & in[455]; 
    assign layer_0[1263] = ~(in[335] ^ in[69]); 
    assign layer_0[1264] = in[395] ^ in[579]; 
    assign layer_0[1265] = ~in[450] | (in[17] & in[450]); 
    assign layer_0[1266] = in[214] ^ in[697]; 
    assign layer_0[1267] = in[534] ^ in[34]; 
    assign layer_0[1268] = ~(in[553] ^ in[710]); 
    assign layer_0[1269] = in[376] & ~in[632]; 
    assign layer_0[1270] = ~in[550]; 
    assign layer_0[1271] = ~in[416] | (in[600] & in[416]); 
    assign layer_0[1272] = in[619] & ~in[636]; 
    assign layer_0[1273] = ~(in[646] ^ in[106]); 
    assign layer_0[1274] = in[364]; 
    assign layer_0[1275] = in[261] ^ in[12]; 
    assign layer_0[1276] = ~(in[598] ^ in[566]); 
    assign layer_0[1277] = in[12]; 
    assign layer_0[1278] = ~(in[590] | in[626]); 
    assign layer_0[1279] = in[550] ^ in[582]; 
    assign layer_0[1280] = ~in[210] | (in[587] & in[210]); 
    assign layer_0[1281] = in[697] & ~in[476]; 
    assign layer_0[1282] = ~(in[553] ^ in[20]); 
    assign layer_0[1283] = ~(in[397] ^ in[461]); 
    assign layer_0[1284] = ~in[234]; 
    assign layer_0[1285] = in[443] | in[195]; 
    assign layer_0[1286] = in[656] ^ in[369]; 
    assign layer_0[1287] = ~in[372]; 
    assign layer_0[1288] = in[650] | in[14]; 
    assign layer_0[1289] = in[225] ^ in[188]; 
    assign layer_0[1290] = in[645] ^ in[62]; 
    assign layer_0[1291] = in[613] ^ in[329]; 
    assign layer_0[1292] = in[663] ^ in[687]; 
    assign layer_0[1293] = ~(in[21] & in[83]); 
    assign layer_0[1294] = ~(in[368] ^ in[647]); 
    assign layer_0[1295] = in[94] & ~in[274]; 
    assign layer_0[1296] = ~(in[45] & in[404]); 
    assign layer_0[1297] = in[344] & in[393]; 
    assign layer_0[1298] = in[760] ^ in[325]; 
    assign layer_0[1299] = in[581] ^ in[651]; 
    assign layer_0[1300] = ~(in[686] & in[352]); 
    assign layer_0[1301] = in[292] & ~in[531]; 
    assign layer_0[1302] = in[142]; 
    assign layer_0[1303] = ~in[195] | (in[195] & in[190]); 
    assign layer_0[1304] = in[457] & ~in[508]; 
    assign layer_0[1305] = in[130] | in[340]; 
    assign layer_0[1306] = ~(in[538] ^ in[42]); 
    assign layer_0[1307] = ~in[436] | (in[436] & in[376]); 
    assign layer_0[1308] = in[94] & in[201]; 
    assign layer_0[1309] = ~in[508]; 
    assign layer_0[1310] = ~(in[694] ^ in[742]); 
    assign layer_0[1311] = in[316] | in[371]; 
    assign layer_0[1312] = ~(in[325] & in[22]); 
    assign layer_0[1313] = in[372] | in[114]; 
    assign layer_0[1314] = ~in[310] | (in[614] & in[310]); 
    assign layer_0[1315] = ~in[452] | (in[564] & in[452]); 
    assign layer_0[1316] = ~in[489] | (in[554] & in[489]); 
    assign layer_0[1317] = ~(in[162] ^ in[186]); 
    assign layer_0[1318] = in[587] ^ in[649]; 
    assign layer_0[1319] = ~(in[371] ^ in[637]); 
    assign layer_0[1320] = in[628] | in[249]; 
    assign layer_0[1321] = in[458] & ~in[432]; 
    assign layer_0[1322] = in[66] & ~in[532]; 
    assign layer_0[1323] = in[381] & ~in[114]; 
    assign layer_0[1324] = ~(in[696] ^ in[243]); 
    assign layer_0[1325] = in[381]; 
    assign layer_0[1326] = in[496] ^ in[633]; 
    assign layer_0[1327] = ~(in[273] | in[424]); 
    assign layer_0[1328] = ~(in[502] | in[141]); 
    assign layer_0[1329] = ~in[220] | (in[220] & in[752]); 
    assign layer_0[1330] = ~in[568] | (in[599] & in[568]); 
    assign layer_0[1331] = ~in[474]; 
    assign layer_0[1332] = ~in[636] | (in[636] & in[687]); 
    assign layer_0[1333] = ~(in[45] ^ in[551]); 
    assign layer_0[1334] = in[342] & in[61]; 
    assign layer_0[1335] = in[85] & ~in[46]; 
    assign layer_0[1336] = ~(in[131] & in[388]); 
    assign layer_0[1337] = ~(in[204] ^ in[639]); 
    assign layer_0[1338] = in[431] | in[100]; 
    assign layer_0[1339] = ~(in[723] ^ in[556]); 
    assign layer_0[1340] = in[113] ^ in[599]; 
    assign layer_0[1341] = ~in[653]; 
    assign layer_0[1342] = ~in[71] | (in[644] & in[71]); 
    assign layer_0[1343] = in[760] | in[322]; 
    assign layer_0[1344] = in[279] ^ in[597]; 
    assign layer_0[1345] = ~in[277] | (in[683] & in[277]); 
    assign layer_0[1346] = ~(in[731] ^ in[550]); 
    assign layer_0[1347] = ~in[262] | (in[553] & in[262]); 
    assign layer_0[1348] = in[599] ^ in[84]; 
    assign layer_0[1349] = ~(in[350] | in[255]); 
    assign layer_0[1350] = in[285] ^ in[449]; 
    assign layer_0[1351] = in[307] ^ in[211]; 
    assign layer_0[1352] = in[30] | in[651]; 
    assign layer_0[1353] = in[692] ^ in[194]; 
    assign layer_0[1354] = ~(in[567] ^ in[581]); 
    assign layer_0[1355] = in[382] & in[143]; 
    assign layer_0[1356] = in[627] & ~in[220]; 
    assign layer_0[1357] = in[485] & in[697]; 
    assign layer_0[1358] = in[120] & ~in[590]; 
    assign layer_0[1359] = in[617] ^ in[420]; 
    assign layer_0[1360] = in[540] | in[722]; 
    assign layer_0[1361] = ~(in[434] ^ in[81]); 
    assign layer_0[1362] = ~(in[552] ^ in[553]); 
    assign layer_0[1363] = in[702] & ~in[615]; 
    assign layer_0[1364] = in[189] ^ in[274]; 
    assign layer_0[1365] = ~in[362]; 
    assign layer_0[1366] = in[630] ^ in[80]; 
    assign layer_0[1367] = ~in[726] | (in[637] & in[726]); 
    assign layer_0[1368] = ~in[539]; 
    assign layer_0[1369] = ~in[487] | (in[487] & in[493]); 
    assign layer_0[1370] = in[229] & in[13]; 
    assign layer_0[1371] = ~in[366]; 
    assign layer_0[1372] = in[632] ^ in[633]; 
    assign layer_0[1373] = ~(in[385] & in[386]); 
    assign layer_0[1374] = ~(in[302] | in[343]); 
    assign layer_0[1375] = ~(in[606] & in[677]); 
    assign layer_0[1376] = in[9]; 
    assign layer_0[1377] = ~in[646] | (in[646] & in[700]); 
    assign layer_0[1378] = in[535] ^ in[744]; 
    assign layer_0[1379] = ~in[238] | (in[550] & in[238]); 
    assign layer_0[1380] = ~in[132]; 
    assign layer_0[1381] = ~(in[587] | in[600]); 
    assign layer_0[1382] = ~in[629]; 
    assign layer_0[1383] = in[717] & ~in[56]; 
    assign layer_0[1384] = in[518]; 
    assign layer_0[1385] = in[9] & in[412]; 
    assign layer_0[1386] = ~(in[492] ^ in[604]); 
    assign layer_0[1387] = in[758] ^ in[603]; 
    assign layer_0[1388] = ~(in[398] | in[104]); 
    assign layer_0[1389] = in[152] & ~in[311]; 
    assign layer_0[1390] = ~(in[693] ^ in[632]); 
    assign layer_0[1391] = in[746]; 
    assign layer_0[1392] = ~in[72]; 
    assign layer_0[1393] = ~in[301] | (in[301] & in[747]); 
    assign layer_0[1394] = in[636] ^ in[703]; 
    assign layer_0[1395] = ~(in[192] & in[404]); 
    assign layer_0[1396] = ~in[509] | (in[408] & in[509]); 
    assign layer_0[1397] = in[380] | in[492]; 
    assign layer_0[1398] = in[78] & in[219]; 
    assign layer_0[1399] = ~in[581]; 
    assign layer_0[1400] = ~(in[751] | in[155]); 
    assign layer_0[1401] = in[278]; 
    assign layer_0[1402] = ~(in[401] | in[407]); 
    assign layer_0[1403] = in[120] & in[86]; 
    assign layer_0[1404] = in[535] & in[362]; 
    assign layer_0[1405] = in[520] | in[293]; 
    assign layer_0[1406] = ~in[598] | (in[760] & in[598]); 
    assign layer_0[1407] = in[629] & ~in[219]; 
    assign layer_0[1408] = in[654] | in[496]; 
    assign layer_0[1409] = in[733] ^ in[204]; 
    assign layer_0[1410] = in[699] | in[570]; 
    assign layer_0[1411] = in[185]; 
    assign layer_0[1412] = ~(in[623] | in[457]); 
    assign layer_0[1413] = in[554] & ~in[697]; 
    assign layer_0[1414] = ~(in[478] | in[519]); 
    assign layer_0[1415] = ~(in[332] | in[246]); 
    assign layer_0[1416] = ~(in[173] | in[647]); 
    assign layer_0[1417] = ~(in[420] ^ in[456]); 
    assign layer_0[1418] = ~(in[506] ^ in[725]); 
    assign layer_0[1419] = ~(in[645] | in[343]); 
    assign layer_0[1420] = in[641] | in[743]; 
    assign layer_0[1421] = in[492] ^ in[244]; 
    assign layer_0[1422] = in[605] ^ in[63]; 
    assign layer_0[1423] = in[475] & in[723]; 
    assign layer_0[1424] = in[669] & ~in[274]; 
    assign layer_0[1425] = ~(in[20] ^ in[158]); 
    assign layer_0[1426] = in[349] | in[28]; 
    assign layer_0[1427] = ~in[647] | (in[647] & in[50]); 
    assign layer_0[1428] = ~in[474]; 
    assign layer_0[1429] = ~(in[626] ^ in[185]); 
    assign layer_0[1430] = ~in[226]; 
    assign layer_0[1431] = 1'b0; 
    assign layer_0[1432] = ~(in[300] ^ in[729]); 
    assign layer_0[1433] = ~(in[686] ^ in[362]); 
    assign layer_0[1434] = ~in[419] | (in[419] & in[591]); 
    assign layer_0[1435] = ~(in[633] | in[524]); 
    assign layer_0[1436] = ~(in[683] ^ in[352]); 
    assign layer_0[1437] = in[468] & ~in[29]; 
    assign layer_0[1438] = ~(in[332] & in[667]); 
    assign layer_0[1439] = ~(in[419] | in[576]); 
    assign layer_0[1440] = ~(in[359] ^ in[266]); 
    assign layer_0[1441] = in[713] ^ in[712]; 
    assign layer_0[1442] = in[578] | in[5]; 
    assign layer_0[1443] = ~(in[419] ^ in[601]); 
    assign layer_0[1444] = ~in[613]; 
    assign layer_0[1445] = in[183] & ~in[234]; 
    assign layer_0[1446] = in[20] & ~in[30]; 
    assign layer_0[1447] = in[85]; 
    assign layer_0[1448] = ~in[38]; 
    assign layer_0[1449] = ~in[766]; 
    assign layer_0[1450] = ~in[519]; 
    assign layer_0[1451] = in[494] & ~in[608]; 
    assign layer_0[1452] = in[367]; 
    assign layer_0[1453] = ~(in[482] ^ in[601]); 
    assign layer_0[1454] = ~(in[582] ^ in[395]); 
    assign layer_0[1455] = ~(in[692] ^ in[727]); 
    assign layer_0[1456] = in[160] & in[603]; 
    assign layer_0[1457] = in[519] | in[667]; 
    assign layer_0[1458] = in[19]; 
    assign layer_0[1459] = in[743]; 
    assign layer_0[1460] = ~(in[92] & in[388]); 
    assign layer_0[1461] = in[736] & ~in[437]; 
    assign layer_0[1462] = in[77] | in[352]; 
    assign layer_0[1463] = ~in[281]; 
    assign layer_0[1464] = in[606] ^ in[434]; 
    assign layer_0[1465] = in[491]; 
    assign layer_0[1466] = in[505] & in[168]; 
    assign layer_0[1467] = in[118] ^ in[196]; 
    assign layer_0[1468] = in[657] & ~in[630]; 
    assign layer_0[1469] = in[662]; 
    assign layer_0[1470] = in[353] ^ in[93]; 
    assign layer_0[1471] = in[1] ^ in[332]; 
    assign layer_0[1472] = in[467] ^ in[212]; 
    assign layer_0[1473] = ~(in[436] ^ in[444]); 
    assign layer_0[1474] = ~(in[583] ^ in[532]); 
    assign layer_0[1475] = ~(in[744] ^ in[646]); 
    assign layer_0[1476] = ~(in[115] & in[599]); 
    assign layer_0[1477] = 1'b0; 
    assign layer_0[1478] = ~(in[484] ^ in[380]); 
    assign layer_0[1479] = in[265] | in[698]; 
    assign layer_0[1480] = ~(in[40] & in[441]); 
    assign layer_0[1481] = in[368] ^ in[746]; 
    assign layer_0[1482] = ~(in[377] & in[582]); 
    assign layer_0[1483] = in[708] & ~in[486]; 
    assign layer_0[1484] = ~(in[473] ^ in[465]); 
    assign layer_0[1485] = ~(in[424] ^ in[286]); 
    assign layer_0[1486] = ~in[650] | (in[650] & in[610]); 
    assign layer_0[1487] = ~(in[122] ^ in[348]); 
    assign layer_0[1488] = in[229] & in[467]; 
    assign layer_0[1489] = in[678]; 
    assign layer_0[1490] = in[401]; 
    assign layer_0[1491] = ~(in[396] & in[407]); 
    assign layer_0[1492] = in[579]; 
    assign layer_0[1493] = ~in[331]; 
    assign layer_0[1494] = in[635] & in[177]; 
    assign layer_0[1495] = ~in[696] | (in[696] & in[161]); 
    assign layer_0[1496] = in[654] & ~in[311]; 
    assign layer_0[1497] = in[620] ^ in[554]; 
    assign layer_0[1498] = ~in[101]; 
    assign layer_0[1499] = ~(in[586] | in[386]); 
    assign layer_0[1500] = ~(in[311] ^ in[580]); 
    assign layer_0[1501] = in[95]; 
    assign layer_0[1502] = in[587] & ~in[312]; 
    assign layer_0[1503] = ~(in[638] & in[653]); 
    assign layer_0[1504] = ~(in[692] ^ in[69]); 
    assign layer_0[1505] = in[612] & in[306]; 
    assign layer_0[1506] = in[673] ^ in[324]; 
    assign layer_0[1507] = ~(in[468] ^ in[483]); 
    assign layer_0[1508] = ~in[382]; 
    assign layer_0[1509] = in[315] & in[691]; 
    assign layer_0[1510] = ~(in[686] ^ in[654]); 
    assign layer_0[1511] = in[537] & ~in[314]; 
    assign layer_0[1512] = in[324]; 
    assign layer_0[1513] = ~(in[33] | in[392]); 
    assign layer_0[1514] = in[407]; 
    assign layer_0[1515] = ~(in[19] ^ in[253]); 
    assign layer_0[1516] = in[695] & ~in[661]; 
    assign layer_0[1517] = ~in[35] | (in[330] & in[35]); 
    assign layer_0[1518] = in[269]; 
    assign layer_0[1519] = ~in[460] | (in[460] & in[740]); 
    assign layer_0[1520] = ~in[335] | (in[600] & in[335]); 
    assign layer_0[1521] = ~in[364]; 
    assign layer_0[1522] = ~in[343] | (in[343] & in[64]); 
    assign layer_0[1523] = in[568] & ~in[655]; 
    assign layer_0[1524] = in[635] & ~in[508]; 
    assign layer_0[1525] = ~in[189] | (in[189] & in[681]); 
    assign layer_0[1526] = ~in[350] | (in[612] & in[350]); 
    assign layer_0[1527] = ~(in[460] & in[396]); 
    assign layer_0[1528] = in[222] | in[401]; 
    assign layer_0[1529] = in[452] | in[618]; 
    assign layer_0[1530] = in[32] | in[502]; 
    assign layer_0[1531] = ~(in[225] ^ in[161]); 
    assign layer_0[1532] = ~in[150] | (in[150] & in[33]); 
    assign layer_0[1533] = in[695] & in[710]; 
    assign layer_0[1534] = in[666]; 
    assign layer_0[1535] = 1'b1; 
    assign layer_0[1536] = in[381]; 
    assign layer_0[1537] = in[230] ^ in[360]; 
    assign layer_0[1538] = in[719] ^ in[99]; 
    assign layer_0[1539] = in[646] & ~in[364]; 
    assign layer_0[1540] = in[60] ^ in[689]; 
    assign layer_0[1541] = ~in[297] | (in[297] & in[650]); 
    assign layer_0[1542] = in[19] & ~in[389]; 
    assign layer_0[1543] = in[709] ^ in[211]; 
    assign layer_0[1544] = ~in[194] | (in[194] & in[261]); 
    assign layer_0[1545] = ~in[379] | (in[647] & in[379]); 
    assign layer_0[1546] = ~(in[45] ^ in[85]); 
    assign layer_0[1547] = in[264] ^ in[604]; 
    assign layer_0[1548] = in[322] ^ in[629]; 
    assign layer_0[1549] = in[377]; 
    assign layer_0[1550] = ~(in[130] & in[316]); 
    assign layer_0[1551] = in[692] ^ in[603]; 
    assign layer_0[1552] = ~(in[197] ^ in[296]); 
    assign layer_0[1553] = ~in[730] | (in[730] & in[98]); 
    assign layer_0[1554] = in[366] & ~in[754]; 
    assign layer_0[1555] = ~(in[615] ^ in[42]); 
    assign layer_0[1556] = ~(in[666] ^ in[645]); 
    assign layer_0[1557] = ~(in[360] & in[636]); 
    assign layer_0[1558] = ~(in[767] | in[659]); 
    assign layer_0[1559] = in[597]; 
    assign layer_0[1560] = 1'b0; 
    assign layer_0[1561] = in[709] & in[296]; 
    assign layer_0[1562] = ~in[554] | (in[18] & in[554]); 
    assign layer_0[1563] = in[217]; 
    assign layer_0[1564] = ~in[12] | (in[12] & in[758]); 
    assign layer_0[1565] = ~(in[220] ^ in[599]); 
    assign layer_0[1566] = ~(in[636] ^ in[177]); 
    assign layer_0[1567] = in[485] ^ in[235]; 
    assign layer_0[1568] = ~in[22] | (in[22] & in[393]); 
    assign layer_0[1569] = ~(in[582] | in[518]); 
    assign layer_0[1570] = ~in[78]; 
    assign layer_0[1571] = ~(in[380] ^ in[109]); 
    assign layer_0[1572] = ~in[321]; 
    assign layer_0[1573] = ~in[569]; 
    assign layer_0[1574] = in[319] ^ in[586]; 
    assign layer_0[1575] = in[205] ^ in[239]; 
    assign layer_0[1576] = ~in[287] | (in[287] & in[90]); 
    assign layer_0[1577] = in[463] ^ in[284]; 
    assign layer_0[1578] = in[187] & ~in[312]; 
    assign layer_0[1579] = in[492] & ~in[47]; 
    assign layer_0[1580] = in[322]; 
    assign layer_0[1581] = in[392]; 
    assign layer_0[1582] = ~in[694]; 
    assign layer_0[1583] = in[200] ^ in[707]; 
    assign layer_0[1584] = ~(in[579] ^ in[475]); 
    assign layer_0[1585] = in[224]; 
    assign layer_0[1586] = ~(in[436] & in[71]); 
    assign layer_0[1587] = ~in[577] | (in[577] & in[165]); 
    assign layer_0[1588] = in[276] & ~in[276]; 
    assign layer_0[1589] = in[643] ^ in[673]; 
    assign layer_0[1590] = ~in[553] | (in[553] & in[300]); 
    assign layer_0[1591] = ~(in[366] | in[641]); 
    assign layer_0[1592] = ~(in[287] | in[156]); 
    assign layer_0[1593] = 1'b0; 
    assign layer_0[1594] = ~in[467] | (in[337] & in[467]); 
    assign layer_0[1595] = ~in[761]; 
    assign layer_0[1596] = ~in[6]; 
    assign layer_0[1597] = ~in[162] | (in[359] & in[162]); 
    assign layer_0[1598] = ~(in[35] | in[19]); 
    assign layer_0[1599] = ~in[399] | (in[629] & in[399]); 
    assign layer_0[1600] = in[692] & ~in[465]; 
    assign layer_0[1601] = in[322] | in[156]; 
    assign layer_0[1602] = in[308] ^ in[412]; 
    assign layer_0[1603] = in[140] ^ in[236]; 
    assign layer_0[1604] = ~(in[142] | in[487]); 
    assign layer_0[1605] = in[206] ^ in[19]; 
    assign layer_0[1606] = ~(in[85] | in[209]); 
    assign layer_0[1607] = ~(in[556] ^ in[546]); 
    assign layer_0[1608] = in[249] & in[489]; 
    assign layer_0[1609] = in[223] ^ in[437]; 
    assign layer_0[1610] = ~(in[3] ^ in[505]); 
    assign layer_0[1611] = in[646] ^ in[719]; 
    assign layer_0[1612] = in[653]; 
    assign layer_0[1613] = in[204]; 
    assign layer_0[1614] = ~in[242] | (in[242] & in[292]); 
    assign layer_0[1615] = in[313] ^ in[291]; 
    assign layer_0[1616] = in[29] | in[312]; 
    assign layer_0[1617] = in[504] ^ in[645]; 
    assign layer_0[1618] = ~in[39] | (in[521] & in[39]); 
    assign layer_0[1619] = in[456] & ~in[207]; 
    assign layer_0[1620] = ~in[644]; 
    assign layer_0[1621] = in[281] ^ in[693]; 
    assign layer_0[1622] = in[384] & ~in[619]; 
    assign layer_0[1623] = ~(in[583] | in[677]); 
    assign layer_0[1624] = in[621] | in[539]; 
    assign layer_0[1625] = in[389] ^ in[315]; 
    assign layer_0[1626] = in[3] ^ in[62]; 
    assign layer_0[1627] = in[149]; 
    assign layer_0[1628] = in[664] ^ in[615]; 
    assign layer_0[1629] = ~(in[404] | in[223]); 
    assign layer_0[1630] = ~(in[51] ^ in[632]); 
    assign layer_0[1631] = ~(in[236] ^ in[600]); 
    assign layer_0[1632] = ~in[316] | (in[316] & in[583]); 
    assign layer_0[1633] = ~in[506] | (in[506] & in[368]); 
    assign layer_0[1634] = ~in[707]; 
    assign layer_0[1635] = ~(in[665] ^ in[580]); 
    assign layer_0[1636] = ~(in[710] ^ in[711]); 
    assign layer_0[1637] = ~in[614]; 
    assign layer_0[1638] = ~(in[39] ^ in[438]); 
    assign layer_0[1639] = in[116]; 
    assign layer_0[1640] = in[670] ^ in[265]; 
    assign layer_0[1641] = ~in[339]; 
    assign layer_0[1642] = in[78] | in[735]; 
    assign layer_0[1643] = in[303]; 
    assign layer_0[1644] = ~in[115] | (in[5] & in[115]); 
    assign layer_0[1645] = in[100] ^ in[693]; 
    assign layer_0[1646] = in[597] & ~in[758]; 
    assign layer_0[1647] = ~in[451] | (in[126] & in[451]); 
    assign layer_0[1648] = in[581] & ~in[594]; 
    assign layer_0[1649] = in[404] ^ in[203]; 
    assign layer_0[1650] = in[78] & ~in[647]; 
    assign layer_0[1651] = ~(in[558] ^ in[69]); 
    assign layer_0[1652] = ~in[497]; 
    assign layer_0[1653] = ~in[473] | (in[473] & in[253]); 
    assign layer_0[1654] = in[617] ^ in[371]; 
    assign layer_0[1655] = in[701] | in[664]; 
    assign layer_0[1656] = ~(in[62] ^ in[476]); 
    assign layer_0[1657] = ~(in[334] ^ in[507]); 
    assign layer_0[1658] = in[600] ^ in[759]; 
    assign layer_0[1659] = in[738]; 
    assign layer_0[1660] = ~in[460]; 
    assign layer_0[1661] = in[375]; 
    assign layer_0[1662] = in[206] ^ in[246]; 
    assign layer_0[1663] = in[571] | in[473]; 
    assign layer_0[1664] = in[581] | in[311]; 
    assign layer_0[1665] = ~in[340]; 
    assign layer_0[1666] = ~(in[276] | in[582]); 
    assign layer_0[1667] = ~in[565]; 
    assign layer_0[1668] = in[311] | in[316]; 
    assign layer_0[1669] = ~in[141] | (in[625] & in[141]); 
    assign layer_0[1670] = in[687]; 
    assign layer_0[1671] = in[595] ^ in[450]; 
    assign layer_0[1672] = ~in[488]; 
    assign layer_0[1673] = ~in[695] | (in[695] & in[45]); 
    assign layer_0[1674] = in[93] ^ in[210]; 
    assign layer_0[1675] = in[652] & ~in[635]; 
    assign layer_0[1676] = ~in[756] | (in[478] & in[756]); 
    assign layer_0[1677] = in[244] & in[299]; 
    assign layer_0[1678] = ~(in[217] | in[507]); 
    assign layer_0[1679] = in[727] & ~in[484]; 
    assign layer_0[1680] = in[633] & ~in[282]; 
    assign layer_0[1681] = ~in[669]; 
    assign layer_0[1682] = ~(in[536] & in[265]); 
    assign layer_0[1683] = ~(in[474] ^ in[581]); 
    assign layer_0[1684] = in[347]; 
    assign layer_0[1685] = in[519] ^ in[315]; 
    assign layer_0[1686] = ~(in[729] ^ in[564]); 
    assign layer_0[1687] = ~(in[583] ^ in[261]); 
    assign layer_0[1688] = in[693] ^ in[427]; 
    assign layer_0[1689] = in[692]; 
    assign layer_0[1690] = in[620] ^ in[655]; 
    assign layer_0[1691] = in[152] | in[562]; 
    assign layer_0[1692] = ~(in[12] ^ in[497]); 
    assign layer_0[1693] = ~(in[472] ^ in[326]); 
    assign layer_0[1694] = ~(in[387] ^ in[581]); 
    assign layer_0[1695] = in[331] ^ in[466]; 
    assign layer_0[1696] = ~in[584] | (in[584] & in[631]); 
    assign layer_0[1697] = in[279]; 
    assign layer_0[1698] = ~in[643] | (in[643] & in[609]); 
    assign layer_0[1699] = in[630] ^ in[330]; 
    assign layer_0[1700] = ~in[7]; 
    assign layer_0[1701] = in[211]; 
    assign layer_0[1702] = in[537] ^ in[60]; 
    assign layer_0[1703] = ~in[45] | (in[45] & in[452]); 
    assign layer_0[1704] = ~(in[661] ^ in[469]); 
    assign layer_0[1705] = in[130] ^ in[192]; 
    assign layer_0[1706] = in[550] ^ in[155]; 
    assign layer_0[1707] = ~(in[372] ^ in[202]); 
    assign layer_0[1708] = ~in[40]; 
    assign layer_0[1709] = in[612]; 
    assign layer_0[1710] = ~in[314] | (in[572] & in[314]); 
    assign layer_0[1711] = ~in[110]; 
    assign layer_0[1712] = in[333] | in[715]; 
    assign layer_0[1713] = ~(in[221] & in[302]); 
    assign layer_0[1714] = in[373]; 
    assign layer_0[1715] = in[28]; 
    assign layer_0[1716] = in[548]; 
    assign layer_0[1717] = ~in[550] | (in[550] & in[284]); 
    assign layer_0[1718] = ~(in[721] ^ in[470]); 
    assign layer_0[1719] = ~(in[237] ^ in[423]); 
    assign layer_0[1720] = in[711] ^ in[335]; 
    assign layer_0[1721] = ~(in[530] | in[365]); 
    assign layer_0[1722] = in[664] & in[300]; 
    assign layer_0[1723] = in[471] | in[184]; 
    assign layer_0[1724] = 1'b1; 
    assign layer_0[1725] = in[415] | in[542]; 
    assign layer_0[1726] = ~(in[243] ^ in[647]); 
    assign layer_0[1727] = in[145] & ~in[569]; 
    assign layer_0[1728] = ~(in[277] ^ in[238]); 
    assign layer_0[1729] = in[344] & in[565]; 
    assign layer_0[1730] = ~(in[316] ^ in[745]); 
    assign layer_0[1731] = in[331] | in[129]; 
    assign layer_0[1732] = in[536]; 
    assign layer_0[1733] = in[407] ^ in[208]; 
    assign layer_0[1734] = ~(in[161] ^ in[190]); 
    assign layer_0[1735] = ~(in[506] ^ in[501]); 
    assign layer_0[1736] = in[598] ^ in[619]; 
    assign layer_0[1737] = in[679] ^ in[273]; 
    assign layer_0[1738] = ~(in[509] ^ in[23]); 
    assign layer_0[1739] = in[45] | in[571]; 
    assign layer_0[1740] = ~(in[332] & in[386]); 
    assign layer_0[1741] = in[226] ^ in[552]; 
    assign layer_0[1742] = in[658]; 
    assign layer_0[1743] = ~in[342] | (in[631] & in[342]); 
    assign layer_0[1744] = in[636] | in[348]; 
    assign layer_0[1745] = ~in[675] | (in[675] & in[10]); 
    assign layer_0[1746] = ~(in[182] & in[300]); 
    assign layer_0[1747] = in[327]; 
    assign layer_0[1748] = ~(in[535] ^ in[170]); 
    assign layer_0[1749] = ~in[387] | (in[254] & in[387]); 
    assign layer_0[1750] = in[316] & in[56]; 
    assign layer_0[1751] = ~(in[710] ^ in[377]); 
    assign layer_0[1752] = ~(in[312] ^ in[657]); 
    assign layer_0[1753] = in[187] | in[459]; 
    assign layer_0[1754] = ~in[597]; 
    assign layer_0[1755] = in[597]; 
    assign layer_0[1756] = in[423] ^ in[384]; 
    assign layer_0[1757] = in[521] & ~in[552]; 
    assign layer_0[1758] = in[316] ^ in[671]; 
    assign layer_0[1759] = in[765]; 
    assign layer_0[1760] = ~(in[12] | in[601]); 
    assign layer_0[1761] = ~(in[262] ^ in[730]); 
    assign layer_0[1762] = in[3] ^ in[628]; 
    assign layer_0[1763] = ~(in[221] & in[331]); 
    assign layer_0[1764] = ~in[631]; 
    assign layer_0[1765] = in[313] ^ in[332]; 
    assign layer_0[1766] = ~(in[731] | in[114]); 
    assign layer_0[1767] = in[145] & in[648]; 
    assign layer_0[1768] = in[146] & ~in[440]; 
    assign layer_0[1769] = in[565]; 
    assign layer_0[1770] = in[339] ^ in[25]; 
    assign layer_0[1771] = ~in[307] | (in[495] & in[307]); 
    assign layer_0[1772] = ~in[596]; 
    assign layer_0[1773] = in[263] ^ in[484]; 
    assign layer_0[1774] = ~(in[615] ^ in[396]); 
    assign layer_0[1775] = ~(in[604] | in[536]); 
    assign layer_0[1776] = in[616]; 
    assign layer_0[1777] = in[685]; 
    assign layer_0[1778] = ~(in[476] & in[617]); 
    assign layer_0[1779] = in[598]; 
    assign layer_0[1780] = ~in[652]; 
    assign layer_0[1781] = in[697] ^ in[555]; 
    assign layer_0[1782] = ~in[645]; 
    assign layer_0[1783] = ~in[307]; 
    assign layer_0[1784] = ~(in[595] ^ in[698]); 
    assign layer_0[1785] = in[426] & ~in[756]; 
    assign layer_0[1786] = ~in[759] | (in[300] & in[759]); 
    assign layer_0[1787] = in[27] & ~in[509]; 
    assign layer_0[1788] = in[725] & ~in[300]; 
    assign layer_0[1789] = in[299] & ~in[263]; 
    assign layer_0[1790] = in[686] & ~in[747]; 
    assign layer_0[1791] = ~(in[411] | in[112]); 
    assign layer_0[1792] = ~in[276] | (in[599] & in[276]); 
    assign layer_0[1793] = in[504]; 
    assign layer_0[1794] = ~(in[533] ^ in[634]); 
    assign layer_0[1795] = ~(in[306] | in[466]); 
    assign layer_0[1796] = in[712] ^ in[430]; 
    assign layer_0[1797] = in[72] & ~in[127]; 
    assign layer_0[1798] = in[732] ^ in[50]; 
    assign layer_0[1799] = ~(in[115] ^ in[145]); 
    assign layer_0[1800] = in[476] & in[619]; 
    assign layer_0[1801] = ~in[744]; 
    assign layer_0[1802] = ~in[38]; 
    assign layer_0[1803] = in[261] & ~in[582]; 
    assign layer_0[1804] = in[550] & ~in[76]; 
    assign layer_0[1805] = in[4] ^ in[507]; 
    assign layer_0[1806] = ~(in[282] ^ in[51]); 
    assign layer_0[1807] = ~(in[487] | in[692]); 
    assign layer_0[1808] = in[328] ^ in[65]; 
    assign layer_0[1809] = in[55]; 
    assign layer_0[1810] = ~in[336]; 
    assign layer_0[1811] = ~(in[450] & in[281]); 
    assign layer_0[1812] = in[761] ^ in[716]; 
    assign layer_0[1813] = in[616] & in[673]; 
    assign layer_0[1814] = in[747]; 
    assign layer_0[1815] = ~(in[291] ^ in[355]); 
    assign layer_0[1816] = ~(in[594] ^ in[247]); 
    assign layer_0[1817] = in[360]; 
    assign layer_0[1818] = ~(in[636] ^ in[430]); 
    assign layer_0[1819] = in[613] & ~in[266]; 
    assign layer_0[1820] = in[166] & in[119]; 
    assign layer_0[1821] = ~(in[174] ^ in[356]); 
    assign layer_0[1822] = in[468] & ~in[762]; 
    assign layer_0[1823] = in[363] & ~in[498]; 
    assign layer_0[1824] = ~(in[158] ^ in[500]); 
    assign layer_0[1825] = ~in[8] | (in[8] & in[762]); 
    assign layer_0[1826] = in[675] ^ in[516]; 
    assign layer_0[1827] = in[443] ^ in[316]; 
    assign layer_0[1828] = ~(in[622] ^ in[638]); 
    assign layer_0[1829] = ~(in[612] ^ in[646]); 
    assign layer_0[1830] = ~(in[478] ^ in[70]); 
    assign layer_0[1831] = ~in[500] | (in[331] & in[500]); 
    assign layer_0[1832] = in[657] ^ in[262]; 
    assign layer_0[1833] = ~(in[395] ^ in[403]); 
    assign layer_0[1834] = in[582]; 
    assign layer_0[1835] = in[634] & ~in[417]; 
    assign layer_0[1836] = in[553] & ~in[368]; 
    assign layer_0[1837] = in[716] & in[409]; 
    assign layer_0[1838] = ~in[536] | (in[584] & in[536]); 
    assign layer_0[1839] = in[289] ^ in[411]; 
    assign layer_0[1840] = in[518]; 
    assign layer_0[1841] = in[235] & ~in[598]; 
    assign layer_0[1842] = ~(in[62] ^ in[418]); 
    assign layer_0[1843] = ~in[577]; 
    assign layer_0[1844] = ~in[29] | (in[428] & in[29]); 
    assign layer_0[1845] = ~in[87] | (in[36] & in[87]); 
    assign layer_0[1846] = ~(in[180] | in[502]); 
    assign layer_0[1847] = in[371] & in[500]; 
    assign layer_0[1848] = ~in[665]; 
    assign layer_0[1849] = in[189]; 
    assign layer_0[1850] = in[4] | in[552]; 
    assign layer_0[1851] = ~in[714]; 
    assign layer_0[1852] = in[582] ^ in[494]; 
    assign layer_0[1853] = in[500] ^ in[260]; 
    assign layer_0[1854] = in[65] ^ in[588]; 
    assign layer_0[1855] = ~(in[600] ^ in[602]); 
    assign layer_0[1856] = ~in[28] | (in[28] & in[649]); 
    assign layer_0[1857] = ~(in[677] ^ in[726]); 
    assign layer_0[1858] = in[171] & ~in[716]; 
    assign layer_0[1859] = in[759] ^ in[760]; 
    assign layer_0[1860] = in[616] ^ in[476]; 
    assign layer_0[1861] = in[492] ^ in[142]; 
    assign layer_0[1862] = ~(in[63] & in[205]); 
    assign layer_0[1863] = in[739] & ~in[734]; 
    assign layer_0[1864] = 1'b1; 
    assign layer_0[1865] = in[502] | in[719]; 
    assign layer_0[1866] = ~in[167] | (in[727] & in[167]); 
    assign layer_0[1867] = in[506] ^ in[300]; 
    assign layer_0[1868] = ~(in[584] & in[277]); 
    assign layer_0[1869] = in[593] | in[519]; 
    assign layer_0[1870] = ~(in[492] ^ in[279]); 
    assign layer_0[1871] = in[260]; 
    assign layer_0[1872] = ~in[299] | (in[251] & in[299]); 
    assign layer_0[1873] = in[566] & ~in[241]; 
    assign layer_0[1874] = ~in[587]; 
    assign layer_0[1875] = in[58] & ~in[761]; 
    assign layer_0[1876] = ~(in[601] ^ in[193]); 
    assign layer_0[1877] = in[231] & ~in[491]; 
    assign layer_0[1878] = in[653] | in[570]; 
    assign layer_0[1879] = ~in[402] | (in[258] & in[402]); 
    assign layer_0[1880] = in[481] & in[172]; 
    assign layer_0[1881] = ~in[51] | (in[51] & in[2]); 
    assign layer_0[1882] = in[409] & in[433]; 
    assign layer_0[1883] = ~(in[458] ^ in[540]); 
    assign layer_0[1884] = ~in[97]; 
    assign layer_0[1885] = ~in[198] | (in[760] & in[198]); 
    assign layer_0[1886] = ~(in[85] ^ in[165]); 
    assign layer_0[1887] = ~in[440]; 
    assign layer_0[1888] = in[245] & in[397]; 
    assign layer_0[1889] = ~in[54]; 
    assign layer_0[1890] = in[283] & in[120]; 
    assign layer_0[1891] = ~in[129] | (in[129] & in[482]); 
    assign layer_0[1892] = in[52] & ~in[540]; 
    assign layer_0[1893] = in[393]; 
    assign layer_0[1894] = ~(in[402] ^ in[612]); 
    assign layer_0[1895] = ~in[369] | (in[209] & in[369]); 
    assign layer_0[1896] = in[665] | in[732]; 
    assign layer_0[1897] = ~(in[94] ^ in[260]); 
    assign layer_0[1898] = ~in[675]; 
    assign layer_0[1899] = ~(in[370] & in[66]); 
    assign layer_0[1900] = ~in[594]; 
    assign layer_0[1901] = in[13] & in[166]; 
    assign layer_0[1902] = in[113] ^ in[582]; 
    assign layer_0[1903] = ~in[418] | (in[273] & in[418]); 
    assign layer_0[1904] = ~in[367] | (in[367] & in[319]); 
    assign layer_0[1905] = in[619] | in[698]; 
    assign layer_0[1906] = in[469] & ~in[547]; 
    assign layer_0[1907] = in[597] ^ in[759]; 
    assign layer_0[1908] = in[62]; 
    assign layer_0[1909] = in[552] ^ in[713]; 
    assign layer_0[1910] = ~(in[250] & in[488]); 
    assign layer_0[1911] = ~in[620] | (in[371] & in[620]); 
    assign layer_0[1912] = in[68]; 
    assign layer_0[1913] = ~(in[204] ^ in[346]); 
    assign layer_0[1914] = ~(in[668] | in[694]); 
    assign layer_0[1915] = ~(in[30] ^ in[338]); 
    assign layer_0[1916] = in[300] ^ in[611]; 
    assign layer_0[1917] = ~in[740] | (in[747] & in[740]); 
    assign layer_0[1918] = in[261] ^ in[364]; 
    assign layer_0[1919] = in[433] ^ in[248]; 
    assign layer_0[1920] = ~(in[714] | in[311]); 
    assign layer_0[1921] = ~in[242] | (in[697] & in[242]); 
    assign layer_0[1922] = ~(in[412] | in[615]); 
    assign layer_0[1923] = in[597] & in[712]; 
    assign layer_0[1924] = in[157] ^ in[533]; 
    assign layer_0[1925] = in[50] ^ in[115]; 
    assign layer_0[1926] = in[507] ^ in[536]; 
    assign layer_0[1927] = ~(in[508] ^ in[228]); 
    assign layer_0[1928] = ~(in[434] ^ in[680]); 
    assign layer_0[1929] = ~in[697]; 
    assign layer_0[1930] = in[697]; 
    assign layer_0[1931] = ~in[418]; 
    assign layer_0[1932] = in[56] ^ in[372]; 
    assign layer_0[1933] = ~(in[555] ^ in[185]); 
    assign layer_0[1934] = ~in[457] | (in[457] & in[507]); 
    assign layer_0[1935] = 1'b0; 
    assign layer_0[1936] = ~(in[690] ^ in[326]); 
    assign layer_0[1937] = in[340] | in[635]; 
    assign layer_0[1938] = ~(in[552] | in[578]); 
    assign layer_0[1939] = ~in[732]; 
    assign layer_0[1940] = ~(in[276] ^ in[667]); 
    assign layer_0[1941] = in[263]; 
    assign layer_0[1942] = ~in[718] | (in[591] & in[718]); 
    assign layer_0[1943] = in[638] & in[59]; 
    assign layer_0[1944] = in[520] ^ in[452]; 
    assign layer_0[1945] = ~(in[651] ^ in[345]); 
    assign layer_0[1946] = ~in[35]; 
    assign layer_0[1947] = in[73] & ~in[152]; 
    assign layer_0[1948] = ~in[683]; 
    assign layer_0[1949] = in[179] & in[5]; 
    assign layer_0[1950] = ~in[176] | (in[604] & in[176]); 
    assign layer_0[1951] = ~in[358]; 
    assign layer_0[1952] = in[485] & ~in[177]; 
    assign layer_0[1953] = ~in[702]; 
    assign layer_0[1954] = ~(in[46] ^ in[651]); 
    assign layer_0[1955] = ~(in[749] ^ in[127]); 
    assign layer_0[1956] = ~in[275]; 
    assign layer_0[1957] = in[328] & ~in[349]; 
    assign layer_0[1958] = ~(in[399] | in[624]); 
    assign layer_0[1959] = ~in[433] | (in[433] & in[719]); 
    assign layer_0[1960] = in[418] ^ in[203]; 
    assign layer_0[1961] = ~(in[547] & in[491]); 
    assign layer_0[1962] = ~in[396]; 
    assign layer_0[1963] = ~(in[618] | in[447]); 
    assign layer_0[1964] = in[322] ^ in[715]; 
    assign layer_0[1965] = in[197] ^ in[40]; 
    assign layer_0[1966] = in[626] & ~in[550]; 
    assign layer_0[1967] = ~(in[549] & in[130]); 
    assign layer_0[1968] = in[746] | in[260]; 
    assign layer_0[1969] = ~(in[238] ^ in[356]); 
    assign layer_0[1970] = ~in[453]; 
    assign layer_0[1971] = ~(in[648] ^ in[71]); 
    assign layer_0[1972] = ~(in[98] ^ in[645]); 
    assign layer_0[1973] = ~in[70] | (in[246] & in[70]); 
    assign layer_0[1974] = ~in[139] | (in[139] & in[68]); 
    assign layer_0[1975] = ~in[594]; 
    assign layer_0[1976] = in[405] & in[194]; 
    assign layer_0[1977] = in[254] ^ in[109]; 
    assign layer_0[1978] = in[509] ^ in[670]; 
    assign layer_0[1979] = in[59] ^ in[603]; 
    assign layer_0[1980] = ~(in[536] ^ in[439]); 
    assign layer_0[1981] = ~in[278]; 
    assign layer_0[1982] = ~(in[5] ^ in[629]); 
    assign layer_0[1983] = ~(in[105] ^ in[60]); 
    assign layer_0[1984] = ~(in[125] ^ in[419]); 
    assign layer_0[1985] = ~(in[203] & in[310]); 
    assign layer_0[1986] = ~(in[628] & in[593]); 
    assign layer_0[1987] = in[115] & ~in[631]; 
    assign layer_0[1988] = ~(in[70] ^ in[5]); 
    assign layer_0[1989] = ~(in[519] ^ in[435]); 
    assign layer_0[1990] = ~in[698]; 
    assign layer_0[1991] = ~(in[599] ^ in[600]); 
    assign layer_0[1992] = ~(in[727] ^ in[292]); 
    assign layer_0[1993] = ~(in[682] | in[276]); 
    assign layer_0[1994] = ~(in[548] & in[254]); 
    assign layer_0[1995] = in[243] | in[744]; 
    assign layer_0[1996] = ~in[645] | (in[645] & in[586]); 
    assign layer_0[1997] = in[468] ^ in[675]; 
    assign layer_0[1998] = ~in[656]; 
    assign layer_0[1999] = ~(in[602] ^ in[619]); 
    assign layer_0[2000] = ~(in[238] & in[238]); 
    assign layer_0[2001] = ~(in[633] ^ in[726]); 
    assign layer_0[2002] = 1'b0; 
    assign layer_0[2003] = in[82] & ~in[196]; 
    assign layer_0[2004] = ~(in[345] ^ in[510]); 
    assign layer_0[2005] = in[9]; 
    assign layer_0[2006] = ~(in[613] & in[483]); 
    assign layer_0[2007] = in[344] & ~in[719]; 
    assign layer_0[2008] = in[387] & ~in[676]; 
    assign layer_0[2009] = ~(in[555] | in[463]); 
    assign layer_0[2010] = ~in[436] | (in[436] & in[759]); 
    assign layer_0[2011] = in[555] & ~in[721]; 
    assign layer_0[2012] = ~in[68]; 
    assign layer_0[2013] = ~(in[472] | in[315]); 
    assign layer_0[2014] = in[458]; 
    assign layer_0[2015] = in[468] | in[538]; 
    assign layer_0[2016] = in[291] ^ in[598]; 
    assign layer_0[2017] = in[140] | in[555]; 
    assign layer_0[2018] = ~(in[251] | in[253]); 
    assign layer_0[2019] = ~in[655] | (in[655] & in[356]); 
    assign layer_0[2020] = in[602] ^ in[509]; 
    assign layer_0[2021] = ~in[395] | (in[395] & in[220]); 
    assign layer_0[2022] = ~in[145]; 
    assign layer_0[2023] = in[684] & in[746]; 
    assign layer_0[2024] = ~(in[692] | in[500]); 
    assign layer_0[2025] = ~in[631] | (in[631] & in[574]); 
    assign layer_0[2026] = in[654] | in[340]; 
    assign layer_0[2027] = in[194]; 
    assign layer_0[2028] = ~(in[518] ^ in[491]); 
    assign layer_0[2029] = in[146]; 
    assign layer_0[2030] = ~(in[342] ^ in[245]); 
    assign layer_0[2031] = ~(in[682] ^ in[666]); 
    assign layer_0[2032] = in[730] ^ in[412]; 
    assign layer_0[2033] = ~in[612]; 
    assign layer_0[2034] = ~in[660]; 
    assign layer_0[2035] = ~(in[262] ^ in[607]); 
    assign layer_0[2036] = ~(in[520] | in[585]); 
    assign layer_0[2037] = in[251] ^ in[759]; 
    assign layer_0[2038] = ~(in[617] ^ in[633]); 
    assign layer_0[2039] = ~in[730]; 
    assign layer_0[2040] = in[0]; 
    assign layer_0[2041] = ~(in[300] ^ in[324]); 
    assign layer_0[2042] = in[248] | in[620]; 
    assign layer_0[2043] = in[361] & ~in[291]; 
    assign layer_0[2044] = 1'b1; 
    assign layer_0[2045] = ~in[743]; 
    assign layer_0[2046] = ~in[547] | (in[547] & in[225]); 
    assign layer_0[2047] = ~(in[744] & in[552]); 
    assign layer_0[2048] = in[730] | in[718]; 
    assign layer_0[2049] = in[317] & ~in[567]; 
    assign layer_0[2050] = in[403] | in[279]; 
    assign layer_0[2051] = ~in[382] | (in[382] & in[611]); 
    assign layer_0[2052] = in[551] | in[249]; 
    assign layer_0[2053] = in[668]; 
    assign layer_0[2054] = ~in[184]; 
    assign layer_0[2055] = in[535]; 
    assign layer_0[2056] = in[193]; 
    assign layer_0[2057] = ~(in[309] ^ in[353]); 
    assign layer_0[2058] = ~(in[761] ^ in[549]); 
    assign layer_0[2059] = ~in[452] | (in[452] & in[77]); 
    assign layer_0[2060] = in[599] ^ in[550]; 
    assign layer_0[2061] = ~(in[661] ^ in[244]); 
    assign layer_0[2062] = in[725] ^ in[726]; 
    assign layer_0[2063] = in[746] ^ in[667]; 
    assign layer_0[2064] = in[380] ^ in[666]; 
    assign layer_0[2065] = in[698] | in[460]; 
    assign layer_0[2066] = in[282] & in[552]; 
    assign layer_0[2067] = ~(in[94] ^ in[44]); 
    assign layer_0[2068] = ~(in[267] & in[437]); 
    assign layer_0[2069] = ~in[618] | (in[611] & in[618]); 
    assign layer_0[2070] = in[715] ^ in[431]; 
    assign layer_0[2071] = ~in[339]; 
    assign layer_0[2072] = ~(in[679] ^ in[536]); 
    assign layer_0[2073] = in[67] | in[15]; 
    assign layer_0[2074] = ~(in[410] & in[690]); 
    assign layer_0[2075] = ~in[113] | (in[113] & in[602]); 
    assign layer_0[2076] = in[232] & ~in[700]; 
    assign layer_0[2077] = in[665] & in[629]; 
    assign layer_0[2078] = in[386] ^ in[352]; 
    assign layer_0[2079] = ~(in[174] & in[353]); 
    assign layer_0[2080] = ~(in[518] | in[622]); 
    assign layer_0[2081] = ~(in[599] ^ in[299]); 
    assign layer_0[2082] = ~in[12]; 
    assign layer_0[2083] = ~(in[352] ^ in[63]); 
    assign layer_0[2084] = ~(in[356] | in[369]); 
    assign layer_0[2085] = ~in[80]; 
    assign layer_0[2086] = ~(in[483] | in[521]); 
    assign layer_0[2087] = ~(in[699] & in[634]); 
    assign layer_0[2088] = in[433] & ~in[640]; 
    assign layer_0[2089] = in[654] & ~in[294]; 
    assign layer_0[2090] = ~(in[585] & in[722]); 
    assign layer_0[2091] = ~(in[760] ^ in[368]); 
    assign layer_0[2092] = ~in[126]; 
    assign layer_0[2093] = in[157] ^ in[650]; 
    assign layer_0[2094] = in[598] | in[431]; 
    assign layer_0[2095] = ~(in[484] | in[90]); 
    assign layer_0[2096] = in[333] | in[63]; 
    assign layer_0[2097] = ~in[539] | (in[539] & in[114]); 
    assign layer_0[2098] = in[618]; 
    assign layer_0[2099] = ~(in[325] & in[626]); 
    assign layer_0[2100] = in[698]; 
    assign layer_0[2101] = in[91] & ~in[253]; 
    assign layer_0[2102] = in[262] | in[60]; 
    assign layer_0[2103] = ~in[643] | (in[643] & in[493]); 
    assign layer_0[2104] = ~in[550]; 
    assign layer_0[2105] = in[742] | in[724]; 
    assign layer_0[2106] = ~in[312] | (in[312] & in[94]); 
    assign layer_0[2107] = ~(in[61] ^ in[161]); 
    assign layer_0[2108] = in[566] | in[342]; 
    assign layer_0[2109] = in[634]; 
    assign layer_0[2110] = ~in[292]; 
    assign layer_0[2111] = ~(in[635] | in[161]); 
    assign layer_0[2112] = in[50] ^ in[551]; 
    assign layer_0[2113] = in[713]; 
    assign layer_0[2114] = ~(in[482] ^ in[618]); 
    assign layer_0[2115] = in[215] & ~in[663]; 
    assign layer_0[2116] = ~(in[639] ^ in[370]); 
    assign layer_0[2117] = in[534] ^ in[539]; 
    assign layer_0[2118] = in[612] ^ in[404]; 
    assign layer_0[2119] = in[611] ^ in[221]; 
    assign layer_0[2120] = ~(in[607] | in[323]); 
    assign layer_0[2121] = in[308] ^ in[708]; 
    assign layer_0[2122] = in[340] & in[279]; 
    assign layer_0[2123] = ~(in[654] ^ in[718]); 
    assign layer_0[2124] = ~(in[385] ^ in[432]); 
    assign layer_0[2125] = in[360] & ~in[334]; 
    assign layer_0[2126] = ~in[756] | (in[756] & in[613]); 
    assign layer_0[2127] = in[387]; 
    assign layer_0[2128] = ~in[739] | (in[681] & in[739]); 
    assign layer_0[2129] = ~(in[557] | in[533]); 
    assign layer_0[2130] = in[326] & ~in[477]; 
    assign layer_0[2131] = in[551] ^ in[420]; 
    assign layer_0[2132] = 1'b1; 
    assign layer_0[2133] = ~(in[308] & in[552]); 
    assign layer_0[2134] = ~(in[743] ^ in[681]); 
    assign layer_0[2135] = in[654]; 
    assign layer_0[2136] = in[709] ^ in[14]; 
    assign layer_0[2137] = in[695] ^ in[322]; 
    assign layer_0[2138] = in[585] & ~in[741]; 
    assign layer_0[2139] = ~in[611]; 
    assign layer_0[2140] = in[169] & ~in[33]; 
    assign layer_0[2141] = in[716] & in[310]; 
    assign layer_0[2142] = ~(in[266] ^ in[338]); 
    assign layer_0[2143] = ~(in[64] | in[396]); 
    assign layer_0[2144] = in[664] | in[10]; 
    assign layer_0[2145] = ~in[304]; 
    assign layer_0[2146] = ~in[630] | (in[221] & in[630]); 
    assign layer_0[2147] = in[582] ^ in[246]; 
    assign layer_0[2148] = in[602]; 
    assign layer_0[2149] = ~in[399] | (in[399] & in[537]); 
    assign layer_0[2150] = ~(in[114] ^ in[740]); 
    assign layer_0[2151] = ~(in[600] & in[534]); 
    assign layer_0[2152] = ~in[116] | (in[116] & in[430]); 
    assign layer_0[2153] = ~in[199] | (in[588] & in[199]); 
    assign layer_0[2154] = ~in[6] | (in[697] & in[6]); 
    assign layer_0[2155] = ~in[343] | (in[520] & in[343]); 
    assign layer_0[2156] = in[604] ^ in[537]; 
    assign layer_0[2157] = ~(in[431] ^ in[214]); 
    assign layer_0[2158] = ~in[434]; 
    assign layer_0[2159] = in[490] ^ in[222]; 
    assign layer_0[2160] = ~(in[474] ^ in[223]); 
    assign layer_0[2161] = ~in[440] | (in[697] & in[440]); 
    assign layer_0[2162] = ~in[333] | (in[239] & in[333]); 
    assign layer_0[2163] = in[95] & in[664]; 
    assign layer_0[2164] = in[720]; 
    assign layer_0[2165] = in[186] & ~in[509]; 
    assign layer_0[2166] = in[366] | in[739]; 
    assign layer_0[2167] = in[40]; 
    assign layer_0[2168] = ~(in[655] ^ in[367]); 
    assign layer_0[2169] = ~(in[201] & in[656]); 
    assign layer_0[2170] = in[692] & ~in[676]; 
    assign layer_0[2171] = ~(in[503] ^ in[115]); 
    assign layer_0[2172] = in[65] ^ in[343]; 
    assign layer_0[2173] = in[265]; 
    assign layer_0[2174] = in[574] | in[512]; 
    assign layer_0[2175] = ~(in[582] ^ in[234]); 
    assign layer_0[2176] = in[726] ^ in[193]; 
    assign layer_0[2177] = ~(in[534] | in[375]); 
    assign layer_0[2178] = in[351] & ~in[602]; 
    assign layer_0[2179] = in[342] & ~in[544]; 
    assign layer_0[2180] = ~in[133] | (in[87] & in[133]); 
    assign layer_0[2181] = ~(in[745] ^ in[744]); 
    assign layer_0[2182] = ~(in[579] | in[510]); 
    assign layer_0[2183] = 1'b0; 
    assign layer_0[2184] = ~(in[645] | in[474]); 
    assign layer_0[2185] = in[188] & ~in[131]; 
    assign layer_0[2186] = in[430] | in[11]; 
    assign layer_0[2187] = ~(in[693] ^ in[491]); 
    assign layer_0[2188] = ~(in[698] & in[332]); 
    assign layer_0[2189] = ~in[650]; 
    assign layer_0[2190] = ~(in[355] | in[681]); 
    assign layer_0[2191] = in[579] & in[265]; 
    assign layer_0[2192] = in[103] & ~in[643]; 
    assign layer_0[2193] = ~(in[211] ^ in[665]); 
    assign layer_0[2194] = in[666] & ~in[372]; 
    assign layer_0[2195] = ~in[158]; 
    assign layer_0[2196] = ~(in[670] ^ in[69]); 
    assign layer_0[2197] = in[332] ^ in[66]; 
    assign layer_0[2198] = ~(in[639] ^ in[671]); 
    assign layer_0[2199] = in[396]; 
    assign layer_0[2200] = in[27] ^ in[69]; 
    assign layer_0[2201] = ~(in[33] & in[397]); 
    assign layer_0[2202] = in[471]; 
    assign layer_0[2203] = ~in[262]; 
    assign layer_0[2204] = ~in[610] | (in[610] & in[601]); 
    assign layer_0[2205] = ~(in[640] ^ in[765]); 
    assign layer_0[2206] = in[602] & ~in[714]; 
    assign layer_0[2207] = in[307] & ~in[450]; 
    assign layer_0[2208] = in[11] | in[596]; 
    assign layer_0[2209] = ~in[66]; 
    assign layer_0[2210] = in[594] ^ in[679]; 
    assign layer_0[2211] = in[333] ^ in[179]; 
    assign layer_0[2212] = ~(in[610] ^ in[628]); 
    assign layer_0[2213] = ~(in[500] | in[351]); 
    assign layer_0[2214] = ~in[389] | (in[389] & in[573]); 
    assign layer_0[2215] = ~(in[507] | in[665]); 
    assign layer_0[2216] = in[23]; 
    assign layer_0[2217] = ~in[441] | (in[441] & in[460]); 
    assign layer_0[2218] = ~in[761]; 
    assign layer_0[2219] = in[567] | in[356]; 
    assign layer_0[2220] = ~in[470]; 
    assign layer_0[2221] = ~(in[277] & in[155]); 
    assign layer_0[2222] = in[216] & ~in[567]; 
    assign layer_0[2223] = ~in[311]; 
    assign layer_0[2224] = ~(in[590] ^ in[192]); 
    assign layer_0[2225] = ~in[326] | (in[326] & in[585]); 
    assign layer_0[2226] = in[45] & ~in[563]; 
    assign layer_0[2227] = in[175] | in[763]; 
    assign layer_0[2228] = in[149] ^ in[174]; 
    assign layer_0[2229] = in[448] & ~in[54]; 
    assign layer_0[2230] = in[411] & ~in[255]; 
    assign layer_0[2231] = in[342] & ~in[530]; 
    assign layer_0[2232] = ~(in[29] ^ in[103]); 
    assign layer_0[2233] = ~in[242] | (in[33] & in[242]); 
    assign layer_0[2234] = ~in[403]; 
    assign layer_0[2235] = ~(in[337] ^ in[493]); 
    assign layer_0[2236] = in[28] ^ in[723]; 
    assign layer_0[2237] = in[714]; 
    assign layer_0[2238] = ~(in[54] ^ in[329]); 
    assign layer_0[2239] = in[665] ^ in[663]; 
    assign layer_0[2240] = in[489] & ~in[461]; 
    assign layer_0[2241] = in[126]; 
    assign layer_0[2242] = ~in[568] | (in[190] & in[568]); 
    assign layer_0[2243] = in[637] & ~in[664]; 
    assign layer_0[2244] = in[248] | in[550]; 
    assign layer_0[2245] = ~(in[292] & in[426]); 
    assign layer_0[2246] = ~(in[5] ^ in[146]); 
    assign layer_0[2247] = in[403]; 
    assign layer_0[2248] = ~in[658] | (in[658] & in[229]); 
    assign layer_0[2249] = ~in[421] | (in[421] & in[2]); 
    assign layer_0[2250] = in[613] ^ in[728]; 
    assign layer_0[2251] = ~(in[730] ^ in[678]); 
    assign layer_0[2252] = ~in[128]; 
    assign layer_0[2253] = in[611] & ~in[417]; 
    assign layer_0[2254] = ~in[355] | (in[625] & in[355]); 
    assign layer_0[2255] = ~(in[303] | in[627]); 
    assign layer_0[2256] = in[440] ^ in[462]; 
    assign layer_0[2257] = in[455] & in[511]; 
    assign layer_0[2258] = ~(in[291] ^ in[230]); 
    assign layer_0[2259] = ~(in[419] ^ in[283]); 
    assign layer_0[2260] = in[147] ^ in[45]; 
    assign layer_0[2261] = in[518] | in[451]; 
    assign layer_0[2262] = ~in[301] | (in[301] & in[267]); 
    assign layer_0[2263] = in[503] ^ in[725]; 
    assign layer_0[2264] = ~(in[725] ^ in[265]); 
    assign layer_0[2265] = in[685] ^ in[458]; 
    assign layer_0[2266] = in[422] & in[360]; 
    assign layer_0[2267] = ~in[732] | (in[732] & in[599]); 
    assign layer_0[2268] = in[104] & ~in[7]; 
    assign layer_0[2269] = in[115] & ~in[487]; 
    assign layer_0[2270] = ~in[22] | (in[22] & in[415]); 
    assign layer_0[2271] = in[146] & ~in[426]; 
    assign layer_0[2272] = in[180] & in[397]; 
    assign layer_0[2273] = ~(in[760] ^ in[294]); 
    assign layer_0[2274] = in[721] ^ in[423]; 
    assign layer_0[2275] = in[567] ^ in[696]; 
    assign layer_0[2276] = ~(in[237] ^ in[46]); 
    assign layer_0[2277] = in[28] ^ in[724]; 
    assign layer_0[2278] = in[317] & ~in[631]; 
    assign layer_0[2279] = ~(in[644] ^ in[673]); 
    assign layer_0[2280] = ~in[291]; 
    assign layer_0[2281] = in[360] & in[328]; 
    assign layer_0[2282] = ~in[50]; 
    assign layer_0[2283] = in[371] & in[292]; 
    assign layer_0[2284] = in[688] | in[750]; 
    assign layer_0[2285] = in[316] & in[382]; 
    assign layer_0[2286] = ~in[34] | (in[34] & in[369]); 
    assign layer_0[2287] = in[663] & ~in[631]; 
    assign layer_0[2288] = in[731] & in[226]; 
    assign layer_0[2289] = in[46] ^ in[36]; 
    assign layer_0[2290] = in[345]; 
    assign layer_0[2291] = ~(in[584] ^ in[583]); 
    assign layer_0[2292] = in[620] | in[496]; 
    assign layer_0[2293] = in[479] ^ in[642]; 
    assign layer_0[2294] = in[22] & in[429]; 
    assign layer_0[2295] = ~(in[689] ^ in[144]); 
    assign layer_0[2296] = in[146]; 
    assign layer_0[2297] = ~(in[725] ^ in[2]); 
    assign layer_0[2298] = in[698] & ~in[68]; 
    assign layer_0[2299] = in[550] & ~in[699]; 
    assign layer_0[2300] = 1'b0; 
    assign layer_0[2301] = ~in[417] | (in[417] & in[644]); 
    assign layer_0[2302] = ~(in[617] ^ in[518]); 
    assign layer_0[2303] = ~in[69]; 
    assign layer_0[2304] = ~(in[388] ^ in[568]); 
    assign layer_0[2305] = ~in[566] | (in[566] & in[292]); 
    assign layer_0[2306] = ~in[79] | (in[79] & in[667]); 
    assign layer_0[2307] = in[619] & in[649]; 
    assign layer_0[2308] = ~in[350] | (in[112] & in[350]); 
    assign layer_0[2309] = in[670] & ~in[311]; 
    assign layer_0[2310] = ~(in[30] ^ in[312]); 
    assign layer_0[2311] = in[326] & ~in[302]; 
    assign layer_0[2312] = in[540] ^ in[611]; 
    assign layer_0[2313] = ~(in[34] ^ in[163]); 
    assign layer_0[2314] = in[94] ^ in[534]; 
    assign layer_0[2315] = in[345] & ~in[318]; 
    assign layer_0[2316] = ~(in[154] | in[582]); 
    assign layer_0[2317] = ~(in[413] ^ in[363]); 
    assign layer_0[2318] = ~(in[551] | in[699]); 
    assign layer_0[2319] = ~(in[169] & in[4]); 
    assign layer_0[2320] = ~in[399] | (in[81] & in[399]); 
    assign layer_0[2321] = in[103] & in[504]; 
    assign layer_0[2322] = in[437]; 
    assign layer_0[2323] = in[318]; 
    assign layer_0[2324] = ~in[372] | (in[713] & in[372]); 
    assign layer_0[2325] = ~(in[611] & in[676]); 
    assign layer_0[2326] = ~in[599] | (in[599] & in[558]); 
    assign layer_0[2327] = ~(in[664] ^ in[666]); 
    assign layer_0[2328] = in[8] | in[661]; 
    assign layer_0[2329] = ~(in[393] & in[13]); 
    assign layer_0[2330] = in[210] & ~in[325]; 
    assign layer_0[2331] = in[582] & in[762]; 
    assign layer_0[2332] = ~(in[341] ^ in[179]); 
    assign layer_0[2333] = in[679] & in[114]; 
    assign layer_0[2334] = in[727] ^ in[758]; 
    assign layer_0[2335] = ~in[613] | (in[497] & in[613]); 
    assign layer_0[2336] = in[745] ^ in[585]; 
    assign layer_0[2337] = in[367] | in[725]; 
    assign layer_0[2338] = in[584] | in[355]; 
    assign layer_0[2339] = ~in[518]; 
    assign layer_0[2340] = ~(in[666] ^ in[81]); 
    assign layer_0[2341] = ~(in[387] | in[462]); 
    assign layer_0[2342] = ~in[86] | (in[528] & in[86]); 
    assign layer_0[2343] = ~in[691]; 
    assign layer_0[2344] = ~in[474] | (in[474] & in[385]); 
    assign layer_0[2345] = in[276]; 
    assign layer_0[2346] = ~(in[393] ^ in[397]); 
    assign layer_0[2347] = ~(in[582] | in[231]); 
    assign layer_0[2348] = in[231]; 
    assign layer_0[2349] = in[427] & in[748]; 
    assign layer_0[2350] = ~in[625]; 
    assign layer_0[2351] = in[712] ^ in[61]; 
    assign layer_0[2352] = in[583] | in[581]; 
    assign layer_0[2353] = in[247] & in[392]; 
    assign layer_0[2354] = ~in[372]; 
    assign layer_0[2355] = in[622] & ~in[537]; 
    assign layer_0[2356] = in[145] ^ in[499]; 
    assign layer_0[2357] = ~in[239]; 
    assign layer_0[2358] = ~(in[328] ^ in[644]); 
    assign layer_0[2359] = ~in[759] | (in[709] & in[759]); 
    assign layer_0[2360] = ~(in[50] ^ in[193]); 
    assign layer_0[2361] = ~in[473] | (in[115] & in[473]); 
    assign layer_0[2362] = in[492] & in[728]; 
    assign layer_0[2363] = ~in[753] | (in[534] & in[753]); 
    assign layer_0[2364] = ~in[698] | (in[519] & in[698]); 
    assign layer_0[2365] = ~(in[364] ^ in[316]); 
    assign layer_0[2366] = in[723]; 
    assign layer_0[2367] = ~(in[282] ^ in[473]); 
    assign layer_0[2368] = ~(in[411] | in[260]); 
    assign layer_0[2369] = ~(in[549] ^ in[502]); 
    assign layer_0[2370] = ~in[703]; 
    assign layer_0[2371] = ~in[707] | (in[98] & in[707]); 
    assign layer_0[2372] = in[142] & ~in[476]; 
    assign layer_0[2373] = in[395] & in[471]; 
    assign layer_0[2374] = ~in[184] | (in[184] & in[670]); 
    assign layer_0[2375] = ~(in[676] ^ in[451]); 
    assign layer_0[2376] = ~(in[696] ^ in[205]); 
    assign layer_0[2377] = ~(in[456] ^ in[406]); 
    assign layer_0[2378] = ~(in[552] ^ in[677]); 
    assign layer_0[2379] = in[652] ^ in[460]; 
    assign layer_0[2380] = in[603] & in[466]; 
    assign layer_0[2381] = ~(in[67] ^ in[620]); 
    assign layer_0[2382] = ~in[760]; 
    assign layer_0[2383] = in[573]; 
    assign layer_0[2384] = in[501]; 
    assign layer_0[2385] = ~in[263]; 
    assign layer_0[2386] = in[418]; 
    assign layer_0[2387] = ~in[609]; 
    assign layer_0[2388] = in[193] & in[210]; 
    assign layer_0[2389] = ~in[424]; 
    assign layer_0[2390] = ~in[647]; 
    assign layer_0[2391] = in[212] ^ in[115]; 
    assign layer_0[2392] = ~in[588]; 
    assign layer_0[2393] = in[714] & in[298]; 
    assign layer_0[2394] = in[357] ^ in[719]; 
    assign layer_0[2395] = ~in[389] | (in[389] & in[603]); 
    assign layer_0[2396] = ~in[38]; 
    assign layer_0[2397] = in[699] ^ in[683]; 
    assign layer_0[2398] = in[460]; 
    assign layer_0[2399] = in[707] ^ in[677]; 
    assign layer_0[2400] = in[619] ^ in[671]; 
    assign layer_0[2401] = in[606] & in[39]; 
    assign layer_0[2402] = ~(in[598] ^ in[341]); 
    assign layer_0[2403] = in[224] & in[235]; 
    assign layer_0[2404] = in[683] | in[419]; 
    assign layer_0[2405] = in[211] & ~in[317]; 
    assign layer_0[2406] = in[8] & in[60]; 
    assign layer_0[2407] = ~in[621] | (in[621] & in[11]); 
    assign layer_0[2408] = in[691] & ~in[699]; 
    assign layer_0[2409] = in[271] & in[303]; 
    assign layer_0[2410] = in[621] & ~in[63]; 
    assign layer_0[2411] = ~(in[638] ^ in[194]); 
    assign layer_0[2412] = in[650] & ~in[618]; 
    assign layer_0[2413] = ~(in[507] ^ in[108]); 
    assign layer_0[2414] = in[474] & ~in[383]; 
    assign layer_0[2415] = in[565] ^ in[346]; 
    assign layer_0[2416] = ~in[74] | (in[443] & in[74]); 
    assign layer_0[2417] = in[522] | in[638]; 
    assign layer_0[2418] = ~in[148]; 
    assign layer_0[2419] = ~in[56] | (in[56] & in[760]); 
    assign layer_0[2420] = ~(in[59] & in[171]); 
    assign layer_0[2421] = in[371] & ~in[729]; 
    assign layer_0[2422] = in[631] ^ in[715]; 
    assign layer_0[2423] = ~(in[223] | in[728]); 
    assign layer_0[2424] = in[720] | in[442]; 
    assign layer_0[2425] = in[698] ^ in[713]; 
    assign layer_0[2426] = in[66]; 
    assign layer_0[2427] = in[74] ^ in[247]; 
    assign layer_0[2428] = in[265] ^ in[713]; 
    assign layer_0[2429] = ~(in[745] ^ in[694]); 
    assign layer_0[2430] = in[75]; 
    assign layer_0[2431] = in[744]; 
    assign layer_0[2432] = in[421] & ~in[446]; 
    assign layer_0[2433] = in[695] ^ in[242]; 
    assign layer_0[2434] = ~(in[112] ^ in[620]); 
    assign layer_0[2435] = ~(in[157] ^ in[326]); 
    assign layer_0[2436] = ~(in[473] & in[474]); 
    assign layer_0[2437] = ~in[617] | (in[57] & in[617]); 
    assign layer_0[2438] = in[712]; 
    assign layer_0[2439] = ~(in[599] | in[467]); 
    assign layer_0[2440] = in[710] & ~in[545]; 
    assign layer_0[2441] = in[333] ^ in[452]; 
    assign layer_0[2442] = ~in[21] | (in[21] & in[467]); 
    assign layer_0[2443] = ~(in[283] & in[410]); 
    assign layer_0[2444] = ~(in[747] ^ in[550]); 
    assign layer_0[2445] = ~(in[478] ^ in[108]); 
    assign layer_0[2446] = ~in[38] | (in[618] & in[38]); 
    assign layer_0[2447] = in[90] & ~in[447]; 
    assign layer_0[2448] = ~(in[30] & in[378]); 
    assign layer_0[2449] = in[744] & in[654]; 
    assign layer_0[2450] = ~in[644] | (in[644] & in[663]); 
    assign layer_0[2451] = ~(in[144] ^ in[465]); 
    assign layer_0[2452] = in[726] | in[347]; 
    assign layer_0[2453] = ~in[61] | (in[267] & in[61]); 
    assign layer_0[2454] = in[457] & in[104]; 
    assign layer_0[2455] = in[189] ^ in[296]; 
    assign layer_0[2456] = in[553]; 
    assign layer_0[2457] = ~in[247]; 
    assign layer_0[2458] = in[389] & in[291]; 
    assign layer_0[2459] = in[441] & ~in[361]; 
    assign layer_0[2460] = ~(in[526] & in[423]); 
    assign layer_0[2461] = in[697]; 
    assign layer_0[2462] = in[708]; 
    assign layer_0[2463] = in[709] & ~in[249]; 
    assign layer_0[2464] = in[100] ^ in[414]; 
    assign layer_0[2465] = ~(in[426] & in[430]); 
    assign layer_0[2466] = ~in[146] | (in[673] & in[146]); 
    assign layer_0[2467] = in[580]; 
    assign layer_0[2468] = ~(in[252] ^ in[676]); 
    assign layer_0[2469] = in[362] | in[545]; 
    assign layer_0[2470] = ~(in[53] ^ in[699]); 
    assign layer_0[2471] = ~in[75]; 
    assign layer_0[2472] = in[14] & ~in[298]; 
    assign layer_0[2473] = in[629] & ~in[59]; 
    assign layer_0[2474] = ~(in[451] & in[279]); 
    assign layer_0[2475] = ~in[329] | (in[329] & in[317]); 
    assign layer_0[2476] = ~(in[680] | in[435]); 
    assign layer_0[2477] = in[322]; 
    assign layer_0[2478] = ~in[291] | (in[291] & in[227]); 
    assign layer_0[2479] = ~(in[284] ^ in[709]); 
    assign layer_0[2480] = in[569]; 
    assign layer_0[2481] = in[639] ^ in[26]; 
    assign layer_0[2482] = in[100]; 
    assign layer_0[2483] = ~in[232] | (in[284] & in[232]); 
    assign layer_0[2484] = ~in[55] | (in[62] & in[55]); 
    assign layer_0[2485] = ~in[679]; 
    assign layer_0[2486] = ~in[508] | (in[110] & in[508]); 
    assign layer_0[2487] = in[714] ^ in[211]; 
    assign layer_0[2488] = ~(in[420] ^ in[443]); 
    assign layer_0[2489] = ~(in[715] ^ in[266]); 
    assign layer_0[2490] = in[359] & ~in[63]; 
    assign layer_0[2491] = ~in[744] | (in[757] & in[744]); 
    assign layer_0[2492] = ~(in[667] & in[243]); 
    assign layer_0[2493] = in[20] & ~in[540]; 
    assign layer_0[2494] = ~(in[683] ^ in[459]); 
    assign layer_0[2495] = ~(in[647] | in[158]); 
    assign layer_0[2496] = in[45] ^ in[644]; 
    assign layer_0[2497] = ~in[521]; 
    assign layer_0[2498] = in[556] & ~in[680]; 
    assign layer_0[2499] = ~(in[293] | in[295]); 
    assign layer_0[2500] = ~(in[646] ^ in[173]); 
    assign layer_0[2501] = in[49] & in[420]; 
    assign layer_0[2502] = ~(in[552] ^ in[645]); 
    assign layer_0[2503] = ~in[617]; 
    assign layer_0[2504] = in[81] & ~in[451]; 
    assign layer_0[2505] = ~(in[456] ^ in[642]); 
    assign layer_0[2506] = ~(in[562] & in[766]); 
    assign layer_0[2507] = in[134] & in[361]; 
    assign layer_0[2508] = in[717] ^ in[162]; 
    assign layer_0[2509] = in[535] ^ in[316]; 
    assign layer_0[2510] = in[59]; 
    assign layer_0[2511] = in[478] & ~in[754]; 
    assign layer_0[2512] = ~(in[34] ^ in[379]); 
    assign layer_0[2513] = ~in[275] | (in[281] & in[275]); 
    assign layer_0[2514] = in[538] ^ in[525]; 
    assign layer_0[2515] = ~(in[276] ^ in[553]); 
    assign layer_0[2516] = ~(in[521] ^ in[609]); 
    assign layer_0[2517] = ~(in[41] ^ in[260]); 
    assign layer_0[2518] = ~in[306]; 
    assign layer_0[2519] = ~(in[235] & in[68]); 
    assign layer_0[2520] = ~in[2] | (in[633] & in[2]); 
    assign layer_0[2521] = in[148] & in[583]; 
    assign layer_0[2522] = in[172] & ~in[38]; 
    assign layer_0[2523] = ~(in[499] | in[44]); 
    assign layer_0[2524] = ~(in[284] | in[716]); 
    assign layer_0[2525] = ~(in[678] ^ in[614]); 
    assign layer_0[2526] = ~(in[705] ^ in[401]); 
    assign layer_0[2527] = in[605] & in[468]; 
    assign layer_0[2528] = ~(in[601] ^ in[312]); 
    assign layer_0[2529] = in[663]; 
    assign layer_0[2530] = in[601] & ~in[215]; 
    assign layer_0[2531] = in[51]; 
    assign layer_0[2532] = ~(in[757] ^ in[638]); 
    assign layer_0[2533] = in[190] & ~in[546]; 
    assign layer_0[2534] = ~in[266]; 
    assign layer_0[2535] = ~in[662] | (in[533] & in[662]); 
    assign layer_0[2536] = in[77] & ~in[267]; 
    assign layer_0[2537] = ~(in[383] & in[234]); 
    assign layer_0[2538] = ~(in[97] | in[177]); 
    assign layer_0[2539] = ~in[215] | (in[215] & in[496]); 
    assign layer_0[2540] = in[213] & ~in[176]; 
    assign layer_0[2541] = in[221] & in[265]; 
    assign layer_0[2542] = in[667] & in[46]; 
    assign layer_0[2543] = in[551] ^ in[604]; 
    assign layer_0[2544] = ~(in[13] | in[94]); 
    assign layer_0[2545] = in[391] | in[114]; 
    assign layer_0[2546] = ~(in[82] & in[567]); 
    assign layer_0[2547] = ~in[468] | (in[447] & in[468]); 
    assign layer_0[2548] = ~(in[102] & in[659]); 
    assign layer_0[2549] = ~in[675] | (in[675] & in[647]); 
    assign layer_0[2550] = in[617] ^ in[531]; 
    assign layer_0[2551] = ~(in[174] ^ in[614]); 
    assign layer_0[2552] = in[178] & ~in[746]; 
    assign layer_0[2553] = ~in[45]; 
    assign layer_0[2554] = in[227] ^ in[292]; 
    assign layer_0[2555] = ~(in[568] & in[694]); 
    assign layer_0[2556] = in[98] | in[745]; 
    assign layer_0[2557] = ~(in[266] ^ in[548]); 
    assign layer_0[2558] = in[676] ^ in[762]; 
    assign layer_0[2559] = ~(in[81] & in[86]); 
    assign layer_0[2560] = in[598] & ~in[601]; 
    assign layer_0[2561] = ~(in[26] ^ in[300]); 
    assign layer_0[2562] = ~in[585] | (in[585] & in[556]); 
    assign layer_0[2563] = in[233] & in[699]; 
    assign layer_0[2564] = ~(in[12] ^ in[222]); 
    assign layer_0[2565] = in[338] & ~in[97]; 
    assign layer_0[2566] = ~(in[615] ^ in[743]); 
    assign layer_0[2567] = ~(in[518] & in[375]); 
    assign layer_0[2568] = ~(in[460] & in[171]); 
    assign layer_0[2569] = in[108] & in[99]; 
    assign layer_0[2570] = 1'b0; 
    assign layer_0[2571] = ~(in[602] ^ in[586]); 
    assign layer_0[2572] = ~in[582] | (in[582] & in[510]); 
    assign layer_0[2573] = ~in[81]; 
    assign layer_0[2574] = in[191] ^ in[327]; 
    assign layer_0[2575] = ~(in[62] | in[506]); 
    assign layer_0[2576] = in[588] | in[596]; 
    assign layer_0[2577] = in[610] ^ in[319]; 
    assign layer_0[2578] = in[239] ^ in[70]; 
    assign layer_0[2579] = in[127]; 
    assign layer_0[2580] = ~(in[172] | in[241]); 
    assign layer_0[2581] = in[422] & ~in[581]; 
    assign layer_0[2582] = in[620] ^ in[740]; 
    assign layer_0[2583] = in[479] ^ in[187]; 
    assign layer_0[2584] = in[402] ^ in[536]; 
    assign layer_0[2585] = in[413] & ~in[3]; 
    assign layer_0[2586] = ~(in[652] | in[637]); 
    assign layer_0[2587] = in[680] | in[760]; 
    assign layer_0[2588] = in[618] & ~in[236]; 
    assign layer_0[2589] = ~(in[343] ^ in[739]); 
    assign layer_0[2590] = in[591] ^ in[277]; 
    assign layer_0[2591] = in[615] | in[689]; 
    assign layer_0[2592] = ~in[104] | (in[104] & in[227]); 
    assign layer_0[2593] = in[614]; 
    assign layer_0[2594] = ~in[631]; 
    assign layer_0[2595] = in[195] & in[593]; 
    assign layer_0[2596] = in[65] | in[324]; 
    assign layer_0[2597] = ~(in[680] | in[265]); 
    assign layer_0[2598] = ~in[451] | (in[451] & in[612]); 
    assign layer_0[2599] = in[400]; 
    assign layer_0[2600] = in[651] & in[612]; 
    assign layer_0[2601] = in[446]; 
    assign layer_0[2602] = in[658] | in[659]; 
    assign layer_0[2603] = in[510] | in[629]; 
    assign layer_0[2604] = in[30]; 
    assign layer_0[2605] = in[665] ^ in[235]; 
    assign layer_0[2606] = in[117] & in[23]; 
    assign layer_0[2607] = ~(in[314] ^ in[669]); 
    assign layer_0[2608] = ~(in[291] ^ in[555]); 
    assign layer_0[2609] = in[233]; 
    assign layer_0[2610] = ~in[379] | (in[94] & in[379]); 
    assign layer_0[2611] = ~in[610]; 
    assign layer_0[2612] = in[264] & ~in[50]; 
    assign layer_0[2613] = in[105] & ~in[630]; 
    assign layer_0[2614] = ~in[39]; 
    assign layer_0[2615] = ~in[15]; 
    assign layer_0[2616] = in[343] ^ in[552]; 
    assign layer_0[2617] = ~(in[570] | in[62]); 
    assign layer_0[2618] = ~(in[727] & in[295]); 
    assign layer_0[2619] = in[410] ^ in[459]; 
    assign layer_0[2620] = in[59] ^ in[517]; 
    assign layer_0[2621] = ~(in[718] ^ in[332]); 
    assign layer_0[2622] = ~(in[135] & in[436]); 
    assign layer_0[2623] = ~(in[392] & in[461]); 
    assign layer_0[2624] = in[145] & in[192]; 
    assign layer_0[2625] = ~(in[355] ^ in[669]); 
    assign layer_0[2626] = ~in[685] | (in[685] & in[524]); 
    assign layer_0[2627] = in[2] ^ in[537]; 
    assign layer_0[2628] = in[630]; 
    assign layer_0[2629] = ~(in[325] & in[618]); 
    assign layer_0[2630] = ~in[72] | (in[192] & in[72]); 
    assign layer_0[2631] = ~(in[15] | in[213]); 
    assign layer_0[2632] = ~(in[674] ^ in[319]); 
    assign layer_0[2633] = ~in[518]; 
    assign layer_0[2634] = ~in[250]; 
    assign layer_0[2635] = ~(in[633] | in[538]); 
    assign layer_0[2636] = ~(in[389] ^ in[295]); 
    assign layer_0[2637] = in[729] ^ in[267]; 
    assign layer_0[2638] = in[110] & ~in[15]; 
    assign layer_0[2639] = in[534] ^ in[412]; 
    assign layer_0[2640] = in[7] | in[613]; 
    assign layer_0[2641] = ~in[37] | (in[37] & in[762]); 
    assign layer_0[2642] = ~(in[534] | in[276]); 
    assign layer_0[2643] = ~(in[190] ^ in[503]); 
    assign layer_0[2644] = in[346]; 
    assign layer_0[2645] = ~in[76] | (in[566] & in[76]); 
    assign layer_0[2646] = ~in[266]; 
    assign layer_0[2647] = ~in[612]; 
    assign layer_0[2648] = ~(in[99] ^ in[364]); 
    assign layer_0[2649] = in[737] | in[613]; 
    assign layer_0[2650] = ~in[218]; 
    assign layer_0[2651] = in[330] ^ in[312]; 
    assign layer_0[2652] = ~(in[3] ^ in[284]); 
    assign layer_0[2653] = in[117] & ~in[68]; 
    assign layer_0[2654] = in[146] & in[417]; 
    assign layer_0[2655] = in[504]; 
    assign layer_0[2656] = in[655] & ~in[672]; 
    assign layer_0[2657] = in[744] & ~in[131]; 
    assign layer_0[2658] = ~(in[698] ^ in[686]); 
    assign layer_0[2659] = ~in[253] | (in[500] & in[253]); 
    assign layer_0[2660] = in[333] | in[560]; 
    assign layer_0[2661] = ~in[491]; 
    assign layer_0[2662] = in[605] & in[702]; 
    assign layer_0[2663] = ~(in[79] & in[72]); 
    assign layer_0[2664] = ~in[105]; 
    assign layer_0[2665] = in[122] ^ in[154]; 
    assign layer_0[2666] = in[255] & ~in[446]; 
    assign layer_0[2667] = ~in[600] | (in[600] & in[31]); 
    assign layer_0[2668] = ~in[400]; 
    assign layer_0[2669] = in[757]; 
    assign layer_0[2670] = ~(in[634] ^ in[668]); 
    assign layer_0[2671] = in[200] & ~in[522]; 
    assign layer_0[2672] = ~in[297] | (in[297] & in[630]); 
    assign layer_0[2673] = ~in[114]; 
    assign layer_0[2674] = in[236] | in[412]; 
    assign layer_0[2675] = in[698] & ~in[640]; 
    assign layer_0[2676] = in[423] & in[167]; 
    assign layer_0[2677] = ~in[340]; 
    assign layer_0[2678] = in[60] | in[535]; 
    assign layer_0[2679] = in[456]; 
    assign layer_0[2680] = ~in[326]; 
    assign layer_0[2681] = ~(in[588] ^ in[713]); 
    assign layer_0[2682] = in[660] & in[408]; 
    assign layer_0[2683] = ~in[424] | (in[424] & in[370]); 
    assign layer_0[2684] = in[483] & ~in[262]; 
    assign layer_0[2685] = ~(in[583] ^ in[710]); 
    assign layer_0[2686] = in[114] ^ in[351]; 
    assign layer_0[2687] = ~(in[114] & in[427]); 
    assign layer_0[2688] = ~in[161] | (in[335] & in[161]); 
    assign layer_0[2689] = ~in[115] | (in[115] & in[729]); 
    assign layer_0[2690] = in[649]; 
    assign layer_0[2691] = ~in[565] | (in[565] & in[672]); 
    assign layer_0[2692] = ~in[160]; 
    assign layer_0[2693] = in[634] ^ in[308]; 
    assign layer_0[2694] = in[616]; 
    assign layer_0[2695] = ~(in[351] ^ in[357]); 
    assign layer_0[2696] = ~(in[172] & in[535]); 
    assign layer_0[2697] = ~(in[564] & in[119]); 
    assign layer_0[2698] = in[657]; 
    assign layer_0[2699] = ~(in[693] ^ in[83]); 
    assign layer_0[2700] = in[164] ^ in[400]; 
    assign layer_0[2701] = ~in[710]; 
    assign layer_0[2702] = in[443] ^ in[632]; 
    assign layer_0[2703] = in[51]; 
    assign layer_0[2704] = in[161] & ~in[501]; 
    assign layer_0[2705] = ~(in[337] | in[350]); 
    assign layer_0[2706] = ~(in[695] ^ in[680]); 
    assign layer_0[2707] = ~in[497] | (in[588] & in[497]); 
    assign layer_0[2708] = in[763] & ~in[626]; 
    assign layer_0[2709] = ~(in[739] ^ in[550]); 
    assign layer_0[2710] = ~in[616]; 
    assign layer_0[2711] = ~in[533]; 
    assign layer_0[2712] = ~(in[423] & in[351]); 
    assign layer_0[2713] = ~in[717] | (in[285] & in[717]); 
    assign layer_0[2714] = in[44] ^ in[715]; 
    assign layer_0[2715] = ~in[82]; 
    assign layer_0[2716] = in[444] ^ in[729]; 
    assign layer_0[2717] = in[95]; 
    assign layer_0[2718] = ~in[428] | (in[428] & in[466]); 
    assign layer_0[2719] = in[619] & ~in[538]; 
    assign layer_0[2720] = ~in[699]; 
    assign layer_0[2721] = in[443] & in[102]; 
    assign layer_0[2722] = ~(in[709] & in[348]); 
    assign layer_0[2723] = in[725]; 
    assign layer_0[2724] = ~(in[217] ^ in[389]); 
    assign layer_0[2725] = ~(in[60] ^ in[268]); 
    assign layer_0[2726] = in[600] ^ in[556]; 
    assign layer_0[2727] = in[321]; 
    assign layer_0[2728] = ~in[678]; 
    assign layer_0[2729] = in[142]; 
    assign layer_0[2730] = in[228] ^ in[638]; 
    assign layer_0[2731] = ~(in[484] | in[159]); 
    assign layer_0[2732] = in[192] ^ in[323]; 
    assign layer_0[2733] = in[249] ^ in[229]; 
    assign layer_0[2734] = ~in[741] | (in[741] & in[564]); 
    assign layer_0[2735] = ~(in[646] ^ in[331]); 
    assign layer_0[2736] = ~(in[744] | in[766]); 
    assign layer_0[2737] = in[112] & ~in[351]; 
    assign layer_0[2738] = 1'b1; 
    assign layer_0[2739] = in[243]; 
    assign layer_0[2740] = ~in[343] | (in[406] & in[343]); 
    assign layer_0[2741] = ~in[379]; 
    assign layer_0[2742] = ~(in[603] ^ in[449]); 
    assign layer_0[2743] = ~(in[50] & in[252]); 
    assign layer_0[2744] = in[100] & ~in[355]; 
    assign layer_0[2745] = ~(in[523] ^ in[444]); 
    assign layer_0[2746] = ~(in[189] ^ in[474]); 
    assign layer_0[2747] = ~in[14]; 
    assign layer_0[2748] = ~(in[727] | in[129]); 
    assign layer_0[2749] = in[647] ^ in[519]; 
    assign layer_0[2750] = ~(in[453] ^ in[238]); 
    assign layer_0[2751] = in[407] & ~in[52]; 
    assign layer_0[2752] = ~in[458]; 
    assign layer_0[2753] = ~in[726]; 
    assign layer_0[2754] = ~in[628]; 
    assign layer_0[2755] = in[99] ^ in[58]; 
    assign layer_0[2756] = in[28] & ~in[284]; 
    assign layer_0[2757] = ~in[301]; 
    assign layer_0[2758] = ~in[621] | (in[766] & in[621]); 
    assign layer_0[2759] = in[367]; 
    assign layer_0[2760] = in[38] & ~in[480]; 
    assign layer_0[2761] = ~in[109] | (in[94] & in[109]); 
    assign layer_0[2762] = ~in[349] | (in[354] & in[349]); 
    assign layer_0[2763] = ~in[695] | (in[695] & in[740]); 
    assign layer_0[2764] = ~(in[393] & in[143]); 
    assign layer_0[2765] = in[57] & in[583]; 
    assign layer_0[2766] = ~(in[182] | in[194]); 
    assign layer_0[2767] = in[539] & ~in[563]; 
    assign layer_0[2768] = in[466] & in[10]; 
    assign layer_0[2769] = ~in[587] | (in[266] & in[587]); 
    assign layer_0[2770] = in[388] & in[162]; 
    assign layer_0[2771] = in[102]; 
    assign layer_0[2772] = in[412] & ~in[755]; 
    assign layer_0[2773] = ~(in[332] ^ in[319]); 
    assign layer_0[2774] = ~(in[488] & in[168]); 
    assign layer_0[2775] = in[394] ^ in[728]; 
    assign layer_0[2776] = in[31] & in[378]; 
    assign layer_0[2777] = in[67] & ~in[389]; 
    assign layer_0[2778] = in[553] & in[266]; 
    assign layer_0[2779] = ~(in[553] ^ in[584]); 
    assign layer_0[2780] = ~in[751]; 
    assign layer_0[2781] = ~(in[77] & in[298]); 
    assign layer_0[2782] = in[23] | in[69]; 
    assign layer_0[2783] = ~in[356]; 
    assign layer_0[2784] = in[665] | in[372]; 
    assign layer_0[2785] = in[714] ^ in[698]; 
    assign layer_0[2786] = ~in[209]; 
    assign layer_0[2787] = ~in[616] | (in[250] & in[616]); 
    assign layer_0[2788] = ~in[580] | (in[274] & in[580]); 
    assign layer_0[2789] = in[571] ^ in[697]; 
    assign layer_0[2790] = ~(in[129] | in[389]); 
    assign layer_0[2791] = ~(in[420] ^ in[45]); 
    assign layer_0[2792] = in[423] & ~in[388]; 
    assign layer_0[2793] = ~(in[140] ^ in[673]); 
    assign layer_0[2794] = in[160]; 
    assign layer_0[2795] = ~in[106]; 
    assign layer_0[2796] = in[296]; 
    assign layer_0[2797] = ~in[744] | (in[717] & in[744]); 
    assign layer_0[2798] = ~(in[567] ^ in[343]); 
    assign layer_0[2799] = ~in[357] | (in[357] & in[582]); 
    assign layer_0[2800] = in[133] & ~in[285]; 
    assign layer_0[2801] = ~(in[757] ^ in[131]); 
    assign layer_0[2802] = ~in[362] | (in[362] & in[584]); 
    assign layer_0[2803] = in[161] & ~in[537]; 
    assign layer_0[2804] = in[580]; 
    assign layer_0[2805] = in[358] & ~in[522]; 
    assign layer_0[2806] = in[596] & ~in[568]; 
    assign layer_0[2807] = ~(in[203] | in[634]); 
    assign layer_0[2808] = in[645] & ~in[18]; 
    assign layer_0[2809] = in[484] ^ in[730]; 
    assign layer_0[2810] = ~(in[407] & in[362]); 
    assign layer_0[2811] = ~(in[66] ^ in[743]); 
    assign layer_0[2812] = ~(in[654] ^ in[24]); 
    assign layer_0[2813] = in[366]; 
    assign layer_0[2814] = ~(in[551] ^ in[387]); 
    assign layer_0[2815] = ~(in[161] | in[145]); 
    assign layer_0[2816] = in[601] & ~in[603]; 
    assign layer_0[2817] = in[215]; 
    assign layer_0[2818] = ~in[417]; 
    assign layer_0[2819] = in[747] ^ in[506]; 
    assign layer_0[2820] = in[119]; 
    assign layer_0[2821] = in[502] ^ in[493]; 
    assign layer_0[2822] = in[87] & ~in[603]; 
    assign layer_0[2823] = in[401] & in[94]; 
    assign layer_0[2824] = in[210] ^ in[370]; 
    assign layer_0[2825] = ~(in[205] ^ in[672]); 
    assign layer_0[2826] = ~(in[639] ^ in[75]); 
    assign layer_0[2827] = ~(in[261] ^ in[436]); 
    assign layer_0[2828] = in[688] | in[83]; 
    assign layer_0[2829] = in[584] ^ in[688]; 
    assign layer_0[2830] = ~in[301] | (in[301] & in[462]); 
    assign layer_0[2831] = ~(in[141] ^ in[460]); 
    assign layer_0[2832] = in[763] | in[638]; 
    assign layer_0[2833] = in[649] & in[637]; 
    assign layer_0[2834] = ~(in[727] ^ in[184]); 
    assign layer_0[2835] = ~(in[283] ^ in[444]); 
    assign layer_0[2836] = 1'b0; 
    assign layer_0[2837] = in[507] ^ in[283]; 
    assign layer_0[2838] = in[205] ^ in[396]; 
    assign layer_0[2839] = in[491] & ~in[334]; 
    assign layer_0[2840] = ~(in[551] ^ in[554]); 
    assign layer_0[2841] = ~(in[120] ^ in[498]); 
    assign layer_0[2842] = in[696] & in[473]; 
    assign layer_0[2843] = ~in[485]; 
    assign layer_0[2844] = in[342] & ~in[350]; 
    assign layer_0[2845] = ~in[661] | (in[661] & in[585]); 
    assign layer_0[2846] = ~in[460] | (in[460] & in[48]); 
    assign layer_0[2847] = ~(in[599] ^ in[567]); 
    assign layer_0[2848] = in[171] & ~in[605]; 
    assign layer_0[2849] = ~(in[473] & in[72]); 
    assign layer_0[2850] = in[656] ^ in[98]; 
    assign layer_0[2851] = ~(in[413] ^ in[80]); 
    assign layer_0[2852] = in[315] ^ in[329]; 
    assign layer_0[2853] = ~in[349]; 
    assign layer_0[2854] = ~in[133]; 
    assign layer_0[2855] = in[135] & ~in[683]; 
    assign layer_0[2856] = ~(in[598] ^ in[585]); 
    assign layer_0[2857] = ~in[582] | (in[582] & in[554]); 
    assign layer_0[2858] = ~in[231] | (in[615] & in[231]); 
    assign layer_0[2859] = ~(in[200] & in[671]); 
    assign layer_0[2860] = ~in[254] | (in[212] & in[254]); 
    assign layer_0[2861] = in[249] ^ in[283]; 
    assign layer_0[2862] = ~in[470] | (in[470] & in[160]); 
    assign layer_0[2863] = ~(in[656] & in[173]); 
    assign layer_0[2864] = ~in[191]; 
    assign layer_0[2865] = ~in[262]; 
    assign layer_0[2866] = ~in[667]; 
    assign layer_0[2867] = in[96] | in[299]; 
    assign layer_0[2868] = ~(in[350] & in[528]); 
    assign layer_0[2869] = in[758]; 
    assign layer_0[2870] = ~(in[733] ^ in[225]); 
    assign layer_0[2871] = in[454] | in[621]; 
    assign layer_0[2872] = in[299]; 
    assign layer_0[2873] = ~in[76] | (in[76] & in[413]); 
    assign layer_0[2874] = in[350] & in[665]; 
    assign layer_0[2875] = in[519] & in[677]; 
    assign layer_0[2876] = ~in[581]; 
    assign layer_0[2877] = ~in[13]; 
    assign layer_0[2878] = ~in[535]; 
    assign layer_0[2879] = 1'b0; 
    assign layer_0[2880] = 1'b0; 
    assign layer_0[2881] = in[457] | in[42]; 
    assign layer_0[2882] = ~(in[670] ^ in[481]); 
    assign layer_0[2883] = ~(in[765] | in[661]); 
    assign layer_0[2884] = in[694] ^ in[671]; 
    assign layer_0[2885] = in[266] | in[522]; 
    assign layer_0[2886] = ~(in[680] ^ in[676]); 
    assign layer_0[2887] = in[752]; 
    assign layer_0[2888] = ~(in[504] & in[334]); 
    assign layer_0[2889] = in[725] ^ in[659]; 
    assign layer_0[2890] = ~(in[537] ^ in[329]); 
    assign layer_0[2891] = ~(in[107] & in[656]); 
    assign layer_0[2892] = in[462] & in[616]; 
    assign layer_0[2893] = ~(in[685] ^ in[473]); 
    assign layer_0[2894] = in[581]; 
    assign layer_0[2895] = in[4]; 
    assign layer_0[2896] = in[640] | in[4]; 
    assign layer_0[2897] = ~in[401] | (in[18] & in[401]); 
    assign layer_0[2898] = in[613] ^ in[618]; 
    assign layer_0[2899] = in[515] & in[556]; 
    assign layer_0[2900] = in[270] ^ in[423]; 
    assign layer_0[2901] = in[498] ^ in[231]; 
    assign layer_0[2902] = in[749] & in[228]; 
    assign layer_0[2903] = ~(in[692] | in[682]); 
    assign layer_0[2904] = in[685] | in[303]; 
    assign layer_0[2905] = in[547]; 
    assign layer_0[2906] = ~(in[697] & in[233]); 
    assign layer_0[2907] = in[331]; 
    assign layer_0[2908] = in[23] ^ in[259]; 
    assign layer_0[2909] = ~in[169] | (in[169] & in[284]); 
    assign layer_0[2910] = ~(in[638] ^ in[54]); 
    assign layer_0[2911] = in[714] ^ in[692]; 
    assign layer_0[2912] = ~(in[92] | in[316]); 
    assign layer_0[2913] = ~(in[575] ^ in[309]); 
    assign layer_0[2914] = ~(in[348] ^ in[636]); 
    assign layer_0[2915] = ~in[312] | (in[312] & in[44]); 
    assign layer_0[2916] = ~(in[695] & in[613]); 
    assign layer_0[2917] = in[260] ^ in[712]; 
    assign layer_0[2918] = in[248] ^ in[675]; 
    assign layer_0[2919] = ~(in[635] | in[724]); 
    assign layer_0[2920] = ~(in[687] | in[42]); 
    assign layer_0[2921] = in[19] & in[190]; 
    assign layer_0[2922] = in[28] | in[188]; 
    assign layer_0[2923] = ~in[351]; 
    assign layer_0[2924] = in[30] & in[207]; 
    assign layer_0[2925] = in[587] | in[387]; 
    assign layer_0[2926] = ~(in[618] | in[628]); 
    assign layer_0[2927] = ~in[25]; 
    assign layer_0[2928] = in[631]; 
    assign layer_0[2929] = ~(in[597] ^ in[521]); 
    assign layer_0[2930] = ~(in[641] ^ in[632]); 
    assign layer_0[2931] = ~in[275]; 
    assign layer_0[2932] = ~in[264] | (in[681] & in[264]); 
    assign layer_0[2933] = ~(in[549] ^ in[659]); 
    assign layer_0[2934] = in[588] ^ in[232]; 
    assign layer_0[2935] = ~(in[518] | in[124]); 
    assign layer_0[2936] = ~(in[28] & in[28]); 
    assign layer_0[2937] = ~in[265]; 
    assign layer_0[2938] = in[652] | in[262]; 
    assign layer_0[2939] = in[277] ^ in[505]; 
    assign layer_0[2940] = in[307] ^ in[619]; 
    assign layer_0[2941] = in[6]; 
    assign layer_0[2942] = in[506] & in[380]; 
    assign layer_0[2943] = ~(in[238] | in[432]); 
    assign layer_0[2944] = ~(in[249] & in[747]); 
    assign layer_0[2945] = ~in[67]; 
    assign layer_0[2946] = ~(in[231] & in[626]); 
    assign layer_0[2947] = ~(in[298] & in[442]); 
    assign layer_0[2948] = in[482] ^ in[603]; 
    assign layer_0[2949] = ~in[51] | (in[320] & in[51]); 
    assign layer_0[2950] = ~(in[588] ^ in[325]); 
    assign layer_0[2951] = ~(in[131] & in[653]); 
    assign layer_0[2952] = in[635]; 
    assign layer_0[2953] = in[661]; 
    assign layer_0[2954] = in[740]; 
    assign layer_0[2955] = ~(in[240] ^ in[226]); 
    assign layer_0[2956] = in[642] ^ in[663]; 
    assign layer_0[2957] = in[58] ^ in[484]; 
    assign layer_0[2958] = ~(in[728] ^ in[208]); 
    assign layer_0[2959] = in[370] | in[434]; 
    assign layer_0[2960] = in[91] & in[460]; 
    assign layer_0[2961] = in[51] & ~in[444]; 
    assign layer_0[2962] = in[362]; 
    assign layer_0[2963] = ~in[596]; 
    assign layer_0[2964] = ~in[552] | (in[552] & in[723]); 
    assign layer_0[2965] = ~in[600] | (in[285] & in[600]); 
    assign layer_0[2966] = ~(in[613] ^ in[250]); 
    assign layer_0[2967] = in[651] ^ in[572]; 
    assign layer_0[2968] = ~(in[470] ^ in[193]); 
    assign layer_0[2969] = ~in[506]; 
    assign layer_0[2970] = in[743]; 
    assign layer_0[2971] = in[324] & ~in[763]; 
    assign layer_0[2972] = in[457] ^ in[600]; 
    assign layer_0[2973] = ~in[595] | (in[595] & in[253]); 
    assign layer_0[2974] = ~in[297]; 
    assign layer_0[2975] = in[637] | in[288]; 
    assign layer_0[2976] = in[447] ^ in[653]; 
    assign layer_0[2977] = ~(in[501] ^ in[110]); 
    assign layer_0[2978] = ~in[265]; 
    assign layer_0[2979] = ~(in[411] | in[648]); 
    assign layer_0[2980] = in[468] ^ in[679]; 
    assign layer_0[2981] = ~(in[589] ^ in[46]); 
    assign layer_0[2982] = in[188] ^ in[589]; 
    assign layer_0[2983] = ~(in[501] ^ in[539]); 
    assign layer_0[2984] = ~in[695]; 
    assign layer_0[2985] = in[483]; 
    assign layer_0[2986] = ~(in[5] ^ in[585]); 
    assign layer_0[2987] = in[653]; 
    assign layer_0[2988] = ~in[302]; 
    assign layer_0[2989] = ~(in[451] | in[291]); 
    assign layer_0[2990] = in[149] & ~in[504]; 
    assign layer_0[2991] = 1'b0; 
    assign layer_0[2992] = ~in[473] | (in[403] & in[473]); 
    assign layer_0[2993] = in[681] ^ in[696]; 
    assign layer_0[2994] = in[476] | in[462]; 
    assign layer_0[2995] = in[696] ^ in[693]; 
    assign layer_0[2996] = in[724]; 
    assign layer_0[2997] = ~(in[389] & in[297]); 
    assign layer_0[2998] = ~(in[238] ^ in[307]); 
    assign layer_0[2999] = ~(in[698] ^ in[652]); 
    assign layer_0[3000] = in[354] ^ in[334]; 
    assign layer_0[3001] = ~(in[67] ^ in[503]); 
    assign layer_0[3002] = ~(in[468] ^ in[85]); 
    assign layer_0[3003] = ~(in[98] | in[539]); 
    assign layer_0[3004] = in[308]; 
    assign layer_0[3005] = ~in[568]; 
    assign layer_0[3006] = ~(in[602] ^ in[599]); 
    assign layer_0[3007] = ~(in[647] ^ in[12]); 
    assign layer_0[3008] = ~in[680] | (in[680] & in[200]); 
    assign layer_0[3009] = in[601] & ~in[8]; 
    assign layer_0[3010] = ~(in[211] | in[763]); 
    assign layer_0[3011] = ~in[698] | (in[698] & in[584]); 
    assign layer_0[3012] = in[499] ^ in[131]; 
    assign layer_0[3013] = ~(in[84] ^ in[726]); 
    assign layer_0[3014] = in[266] ^ in[758]; 
    assign layer_0[3015] = in[727] | in[726]; 
    assign layer_0[3016] = in[150] ^ in[558]; 
    assign layer_0[3017] = ~in[177]; 
    assign layer_0[3018] = 1'b1; 
    assign layer_0[3019] = in[710] & ~in[12]; 
    assign layer_0[3020] = in[605]; 
    assign layer_0[3021] = in[55] ^ in[733]; 
    assign layer_0[3022] = ~(in[158] ^ in[412]); 
    assign layer_0[3023] = in[30] ^ in[43]; 
    assign layer_0[3024] = ~in[331] | (in[722] & in[331]); 
    assign layer_0[3025] = ~in[555]; 
    assign layer_0[3026] = in[535] & ~in[338]; 
    assign layer_0[3027] = 1'b0; 
    assign layer_0[3028] = in[476] & ~in[728]; 
    assign layer_0[3029] = ~(in[10] | in[584]); 
    assign layer_0[3030] = in[233] & ~in[722]; 
    assign layer_0[3031] = in[648] & ~in[630]; 
    assign layer_0[3032] = ~(in[235] ^ in[406]); 
    assign layer_0[3033] = in[630] & ~in[75]; 
    assign layer_0[3034] = in[632] & ~in[751]; 
    assign layer_0[3035] = ~(in[296] & in[82]); 
    assign layer_0[3036] = ~(in[719] & in[190]); 
    assign layer_0[3037] = ~in[212] | (in[212] & in[674]); 
    assign layer_0[3038] = in[632] & ~in[758]; 
    assign layer_0[3039] = ~in[326] | (in[326] & in[765]); 
    assign layer_0[3040] = in[265] ^ in[534]; 
    assign layer_0[3041] = in[390] & ~in[248]; 
    assign layer_0[3042] = ~(in[574] ^ in[723]); 
    assign layer_0[3043] = ~in[489] | (in[489] & in[747]); 
    assign layer_0[3044] = in[316] ^ in[111]; 
    assign layer_0[3045] = ~in[617] | (in[688] & in[617]); 
    assign layer_0[3046] = ~(in[229] | in[656]); 
    assign layer_0[3047] = in[277] & ~in[445]; 
    assign layer_0[3048] = ~(in[405] ^ in[338]); 
    assign layer_0[3049] = ~(in[661] ^ in[603]); 
    assign layer_0[3050] = in[404] ^ in[435]; 
    assign layer_0[3051] = in[520] ^ in[99]; 
    assign layer_0[3052] = ~in[684] | (in[697] & in[684]); 
    assign layer_0[3053] = ~in[746]; 
    assign layer_0[3054] = in[534] | in[625]; 
    assign layer_0[3055] = in[663] & in[404]; 
    assign layer_0[3056] = in[118] | in[727]; 
    assign layer_0[3057] = ~(in[487] & in[627]); 
    assign layer_0[3058] = ~in[634] | (in[372] & in[634]); 
    assign layer_0[3059] = in[699] ^ in[741]; 
    assign layer_0[3060] = ~(in[234] | in[225]); 
    assign layer_0[3061] = in[661] & ~in[221]; 
    assign layer_0[3062] = in[364] & in[404]; 
    assign layer_0[3063] = ~in[451] | (in[451] & in[262]); 
    assign layer_0[3064] = in[263] & in[281]; 
    assign layer_0[3065] = ~(in[661] | in[384]); 
    assign layer_0[3066] = in[493]; 
    assign layer_0[3067] = in[355] ^ in[421]; 
    assign layer_0[3068] = in[316] ^ in[314]; 
    assign layer_0[3069] = in[388]; 
    assign layer_0[3070] = in[385] & ~in[739]; 
    assign layer_0[3071] = ~(in[131] ^ in[178]); 
    assign layer_0[3072] = ~(in[725] & in[501]); 
    assign layer_0[3073] = in[380]; 
    assign layer_0[3074] = in[106] & ~in[219]; 
    assign layer_0[3075] = ~(in[581] & in[744]); 
    assign layer_0[3076] = ~(in[323] & in[50]); 
    assign layer_0[3077] = ~(in[387] ^ in[162]); 
    assign layer_0[3078] = in[602] & ~in[504]; 
    assign layer_0[3079] = in[743] ^ in[742]; 
    assign layer_0[3080] = in[440]; 
    assign layer_0[3081] = ~(in[111] ^ in[762]); 
    assign layer_0[3082] = in[638]; 
    assign layer_0[3083] = in[405] ^ in[13]; 
    assign layer_0[3084] = in[610] ^ in[392]; 
    assign layer_0[3085] = in[46]; 
    assign layer_0[3086] = in[267] ^ in[263]; 
    assign layer_0[3087] = ~(in[367] & in[611]); 
    assign layer_0[3088] = in[173] ^ in[155]; 
    assign layer_0[3089] = in[597] ^ in[322]; 
    assign layer_0[3090] = ~in[186] | (in[186] & in[689]); 
    assign layer_0[3091] = ~(in[632] ^ in[482]); 
    assign layer_0[3092] = in[486] & ~in[193]; 
    assign layer_0[3093] = ~in[30]; 
    assign layer_0[3094] = in[650] & ~in[697]; 
    assign layer_0[3095] = in[690] ^ in[448]; 
    assign layer_0[3096] = in[667] ^ in[696]; 
    assign layer_0[3097] = in[504] ^ in[483]; 
    assign layer_0[3098] = ~in[56] | (in[479] & in[56]); 
    assign layer_0[3099] = in[753] | in[341]; 
    assign layer_0[3100] = ~in[97]; 
    assign layer_0[3101] = ~in[452] | (in[331] & in[452]); 
    assign layer_0[3102] = ~in[7]; 
    assign layer_0[3103] = in[404]; 
    assign layer_0[3104] = in[420] & ~in[493]; 
    assign layer_0[3105] = ~(in[387] | in[459]); 
    assign layer_0[3106] = ~in[110] | (in[532] & in[110]); 
    assign layer_0[3107] = in[476] ^ in[324]; 
    assign layer_0[3108] = ~in[728] | (in[728] & in[74]); 
    assign layer_0[3109] = in[504] ^ in[298]; 
    assign layer_0[3110] = ~(in[669] | in[486]); 
    assign layer_0[3111] = ~(in[538] | in[758]); 
    assign layer_0[3112] = in[98] & ~in[267]; 
    assign layer_0[3113] = in[282] & ~in[681]; 
    assign layer_0[3114] = ~(in[712] ^ in[744]); 
    assign layer_0[3115] = ~in[205] | (in[728] & in[205]); 
    assign layer_0[3116] = in[462] ^ in[351]; 
    assign layer_0[3117] = in[726] & ~in[731]; 
    assign layer_0[3118] = ~(in[460] ^ in[410]); 
    assign layer_0[3119] = ~(in[492] & in[225]); 
    assign layer_0[3120] = ~in[82]; 
    assign layer_0[3121] = in[424] & in[406]; 
    assign layer_0[3122] = in[315] & in[728]; 
    assign layer_0[3123] = in[106] & ~in[373]; 
    assign layer_0[3124] = in[615] | in[3]; 
    assign layer_0[3125] = in[697] & ~in[597]; 
    assign layer_0[3126] = in[404] & ~in[469]; 
    assign layer_0[3127] = in[347] & in[499]; 
    assign layer_0[3128] = in[760] & ~in[285]; 
    assign layer_0[3129] = in[549]; 
    assign layer_0[3130] = ~(in[461] | in[134]); 
    assign layer_0[3131] = ~(in[452] ^ in[174]); 
    assign layer_0[3132] = ~(in[329] ^ in[685]); 
    assign layer_0[3133] = in[159] & in[452]; 
    assign layer_0[3134] = in[140] ^ in[554]; 
    assign layer_0[3135] = in[730] | in[692]; 
    assign layer_0[3136] = in[646] ^ in[615]; 
    assign layer_0[3137] = in[502] ^ in[678]; 
    assign layer_0[3138] = in[755] ^ in[341]; 
    assign layer_0[3139] = ~(in[741] ^ in[159]); 
    assign layer_0[3140] = ~in[471]; 
    assign layer_0[3141] = ~in[208]; 
    assign layer_0[3142] = ~in[441] | (in[441] & in[109]); 
    assign layer_0[3143] = ~in[84]; 
    assign layer_0[3144] = in[533] | in[222]; 
    assign layer_0[3145] = in[331] & ~in[477]; 
    assign layer_0[3146] = ~in[457] | (in[534] & in[457]); 
    assign layer_0[3147] = ~(in[586] ^ in[215]); 
    assign layer_0[3148] = in[233] ^ in[481]; 
    assign layer_0[3149] = ~(in[349] ^ in[81]); 
    assign layer_0[3150] = in[127] ^ in[635]; 
    assign layer_0[3151] = in[5] ^ in[478]; 
    assign layer_0[3152] = ~in[243]; 
    assign layer_0[3153] = ~in[699] | (in[486] & in[699]); 
    assign layer_0[3154] = ~(in[461] ^ in[230]); 
    assign layer_0[3155] = in[403] ^ in[684]; 
    assign layer_0[3156] = in[392] ^ in[372]; 
    assign layer_0[3157] = ~(in[324] ^ in[116]); 
    assign layer_0[3158] = ~(in[681] ^ in[333]); 
    assign layer_0[3159] = in[253] ^ in[475]; 
    assign layer_0[3160] = in[404] ^ in[552]; 
    assign layer_0[3161] = in[254]; 
    assign layer_0[3162] = in[92] & in[124]; 
    assign layer_0[3163] = in[722] ^ in[425]; 
    assign layer_0[3164] = ~in[381] | (in[381] & in[574]); 
    assign layer_0[3165] = ~in[548]; 
    assign layer_0[3166] = ~in[711] | (in[711] & in[530]); 
    assign layer_0[3167] = in[403] & ~in[477]; 
    assign layer_0[3168] = in[650] | in[591]; 
    assign layer_0[3169] = in[693] & in[41]; 
    assign layer_0[3170] = in[51]; 
    assign layer_0[3171] = in[322] ^ in[610]; 
    assign layer_0[3172] = ~(in[634] ^ in[636]); 
    assign layer_0[3173] = in[695] | in[237]; 
    assign layer_0[3174] = in[630] ^ in[663]; 
    assign layer_0[3175] = ~in[708] | (in[708] & in[536]); 
    assign layer_0[3176] = in[604] ^ in[280]; 
    assign layer_0[3177] = ~in[59]; 
    assign layer_0[3178] = in[341]; 
    assign layer_0[3179] = in[365]; 
    assign layer_0[3180] = in[82]; 
    assign layer_0[3181] = in[488] ^ in[28]; 
    assign layer_0[3182] = in[360] & ~in[433]; 
    assign layer_0[3183] = in[301]; 
    assign layer_0[3184] = ~in[441] | (in[441] & in[701]); 
    assign layer_0[3185] = ~(in[744] & in[490]); 
    assign layer_0[3186] = in[644] & ~in[684]; 
    assign layer_0[3187] = ~in[391] | (in[354] & in[391]); 
    assign layer_0[3188] = in[488] & ~in[502]; 
    assign layer_0[3189] = ~(in[492] & in[145]); 
    assign layer_0[3190] = ~in[79] | (in[79] & in[572]); 
    assign layer_0[3191] = in[520] ^ in[762]; 
    assign layer_0[3192] = in[224] ^ in[492]; 
    assign layer_0[3193] = in[568]; 
    assign layer_0[3194] = ~(in[352] | in[605]); 
    assign layer_0[3195] = ~in[666] | (in[301] & in[666]); 
    assign layer_0[3196] = ~(in[162] ^ in[3]); 
    assign layer_0[3197] = ~(in[241] | in[588]); 
    assign layer_0[3198] = in[194] | in[614]; 
    assign layer_0[3199] = in[295] | in[294]; 
    assign layer_0[3200] = ~(in[267] | in[466]); 
    assign layer_0[3201] = ~(in[298] | in[608]); 
    assign layer_0[3202] = in[552] ^ in[550]; 
    assign layer_0[3203] = in[460] ^ in[200]; 
    assign layer_0[3204] = in[662] & in[535]; 
    assign layer_0[3205] = ~(in[292] ^ in[483]); 
    assign layer_0[3206] = ~(in[645] | in[135]); 
    assign layer_0[3207] = ~in[162] | (in[94] & in[162]); 
    assign layer_0[3208] = ~in[570]; 
    assign layer_0[3209] = in[261] | in[458]; 
    assign layer_0[3210] = ~(in[705] ^ in[670]); 
    assign layer_0[3211] = ~in[631]; 
    assign layer_0[3212] = ~(in[424] | in[404]); 
    assign layer_0[3213] = in[538] ^ in[743]; 
    assign layer_0[3214] = in[572] ^ in[365]; 
    assign layer_0[3215] = in[502]; 
    assign layer_0[3216] = ~(in[220] ^ in[253]); 
    assign layer_0[3217] = ~in[354]; 
    assign layer_0[3218] = in[535] ^ in[315]; 
    assign layer_0[3219] = ~(in[20] | in[44]); 
    assign layer_0[3220] = in[451] ^ in[7]; 
    assign layer_0[3221] = in[659] ^ in[313]; 
    assign layer_0[3222] = in[41] & in[18]; 
    assign layer_0[3223] = ~in[61] | (in[61] & in[668]); 
    assign layer_0[3224] = in[483] & in[291]; 
    assign layer_0[3225] = ~(in[727] ^ in[264]); 
    assign layer_0[3226] = ~(in[277] ^ in[760]); 
    assign layer_0[3227] = in[619]; 
    assign layer_0[3228] = in[423] ^ in[588]; 
    assign layer_0[3229] = in[61] & ~in[189]; 
    assign layer_0[3230] = ~in[567] | (in[128] & in[567]); 
    assign layer_0[3231] = ~in[624]; 
    assign layer_0[3232] = ~(in[136] ^ in[144]); 
    assign layer_0[3233] = in[252] ^ in[551]; 
    assign layer_0[3234] = ~(in[250] & in[444]); 
    assign layer_0[3235] = in[614] & ~in[432]; 
    assign layer_0[3236] = ~in[734]; 
    assign layer_0[3237] = ~in[300] | (in[300] & in[710]); 
    assign layer_0[3238] = in[667] ^ in[586]; 
    assign layer_0[3239] = ~in[98]; 
    assign layer_0[3240] = ~(in[500] | in[452]); 
    assign layer_0[3241] = ~(in[708] ^ in[672]); 
    assign layer_0[3242] = ~(in[596] ^ in[339]); 
    assign layer_0[3243] = ~in[282]; 
    assign layer_0[3244] = in[44]; 
    assign layer_0[3245] = ~in[131]; 
    assign layer_0[3246] = in[340]; 
    assign layer_0[3247] = ~in[475] | (in[523] & in[475]); 
    assign layer_0[3248] = in[5] & ~in[191]; 
    assign layer_0[3249] = in[452] ^ in[731]; 
    assign layer_0[3250] = ~in[266] | (in[760] & in[266]); 
    assign layer_0[3251] = in[333] | in[603]; 
    assign layer_0[3252] = ~(in[54] & in[380]); 
    assign layer_0[3253] = ~(in[677] | in[585]); 
    assign layer_0[3254] = ~(in[650] | in[284]); 
    assign layer_0[3255] = in[465]; 
    assign layer_0[3256] = in[347] & ~in[562]; 
    assign layer_0[3257] = ~(in[290] | in[606]); 
    assign layer_0[3258] = in[699] | in[301]; 
    assign layer_0[3259] = ~(in[195] | in[628]); 
    assign layer_0[3260] = in[192]; 
    assign layer_0[3261] = in[514] ^ in[95]; 
    assign layer_0[3262] = ~in[650]; 
    assign layer_0[3263] = in[747] ^ in[146]; 
    assign layer_0[3264] = in[174] & ~in[668]; 
    assign layer_0[3265] = ~(in[712] ^ in[728]); 
    assign layer_0[3266] = in[341] ^ in[129]; 
    assign layer_0[3267] = in[602] & ~in[561]; 
    assign layer_0[3268] = in[348]; 
    assign layer_0[3269] = in[126] ^ in[629]; 
    assign layer_0[3270] = ~in[374] | (in[374] & in[628]); 
    assign layer_0[3271] = ~in[698]; 
    assign layer_0[3272] = in[754] ^ in[626]; 
    assign layer_0[3273] = ~in[3]; 
    assign layer_0[3274] = ~in[470]; 
    assign layer_0[3275] = in[201] & ~in[78]; 
    assign layer_0[3276] = in[327]; 
    assign layer_0[3277] = ~(in[3] & in[198]); 
    assign layer_0[3278] = ~in[67]; 
    assign layer_0[3279] = in[538] ^ in[395]; 
    assign layer_0[3280] = in[187] & in[349]; 
    assign layer_0[3281] = in[3] ^ in[641]; 
    assign layer_0[3282] = ~(in[635] ^ in[652]); 
    assign layer_0[3283] = in[614] ^ in[759]; 
    assign layer_0[3284] = ~(in[679] & in[425]); 
    assign layer_0[3285] = in[92] ^ in[307]; 
    assign layer_0[3286] = in[740] & ~in[337]; 
    assign layer_0[3287] = in[572] & in[611]; 
    assign layer_0[3288] = in[758] ^ in[131]; 
    assign layer_0[3289] = ~(in[356] | in[435]); 
    assign layer_0[3290] = ~(in[157] | in[307]); 
    assign layer_0[3291] = in[115] & ~in[287]; 
    assign layer_0[3292] = ~(in[139] & in[51]); 
    assign layer_0[3293] = in[40] ^ in[177]; 
    assign layer_0[3294] = in[488] ^ in[20]; 
    assign layer_0[3295] = in[210] ^ in[62]; 
    assign layer_0[3296] = ~(in[595] & in[5]); 
    assign layer_0[3297] = ~in[390] | (in[390] & in[502]); 
    assign layer_0[3298] = in[431] & ~in[630]; 
    assign layer_0[3299] = ~in[663] | (in[663] & in[483]); 
    assign layer_0[3300] = ~in[238] | (in[238] & in[726]); 
    assign layer_0[3301] = in[698] ^ in[432]; 
    assign layer_0[3302] = in[620]; 
    assign layer_0[3303] = ~in[392] | (in[531] & in[392]); 
    assign layer_0[3304] = ~(in[161] ^ in[363]); 
    assign layer_0[3305] = in[147] & ~in[448]; 
    assign layer_0[3306] = in[419]; 
    assign layer_0[3307] = in[328] ^ in[79]; 
    assign layer_0[3308] = in[638] ^ in[216]; 
    assign layer_0[3309] = ~(in[740] | in[144]); 
    assign layer_0[3310] = in[25] & ~in[605]; 
    assign layer_0[3311] = in[244] ^ in[482]; 
    assign layer_0[3312] = ~(in[648] ^ in[189]); 
    assign layer_0[3313] = ~in[579] | (in[511] & in[579]); 
    assign layer_0[3314] = ~(in[761] ^ in[757]); 
    assign layer_0[3315] = ~(in[333] | in[468]); 
    assign layer_0[3316] = ~in[650]; 
    assign layer_0[3317] = ~(in[599] ^ in[612]); 
    assign layer_0[3318] = ~in[245] | (in[245] & in[540]); 
    assign layer_0[3319] = in[641] | in[458]; 
    assign layer_0[3320] = in[282] ^ in[600]; 
    assign layer_0[3321] = ~(in[26] & in[123]); 
    assign layer_0[3322] = in[740] ^ in[282]; 
    assign layer_0[3323] = ~(in[23] ^ in[348]); 
    assign layer_0[3324] = ~in[332] | (in[332] & in[729]); 
    assign layer_0[3325] = in[612] | in[339]; 
    assign layer_0[3326] = in[198] ^ in[601]; 
    assign layer_0[3327] = ~in[267] | (in[267] & in[523]); 
    assign layer_0[3328] = in[435] & ~in[339]; 
    assign layer_0[3329] = ~(in[633] ^ in[602]); 
    assign layer_0[3330] = in[223] ^ in[539]; 
    assign layer_0[3331] = ~(in[650] ^ in[251]); 
    assign layer_0[3332] = in[450] & ~in[518]; 
    assign layer_0[3333] = in[676] & in[326]; 
    assign layer_0[3334] = ~in[100]; 
    assign layer_0[3335] = ~(in[692] ^ in[729]); 
    assign layer_0[3336] = 1'b0; 
    assign layer_0[3337] = ~in[38]; 
    assign layer_0[3338] = ~(in[477] ^ in[469]); 
    assign layer_0[3339] = in[446]; 
    assign layer_0[3340] = in[147] ^ in[689]; 
    assign layer_0[3341] = in[279] ^ in[696]; 
    assign layer_0[3342] = in[588] & in[458]; 
    assign layer_0[3343] = in[762] ^ in[533]; 
    assign layer_0[3344] = in[175] | in[223]; 
    assign layer_0[3345] = in[614] & ~in[158]; 
    assign layer_0[3346] = ~in[428]; 
    assign layer_0[3347] = in[760]; 
    assign layer_0[3348] = in[291]; 
    assign layer_0[3349] = in[235] ^ in[568]; 
    assign layer_0[3350] = in[428] | in[428]; 
    assign layer_0[3351] = ~(in[673] ^ in[644]); 
    assign layer_0[3352] = ~(in[396] ^ in[537]); 
    assign layer_0[3353] = in[356] ^ in[415]; 
    assign layer_0[3354] = 1'b1; 
    assign layer_0[3355] = in[333] & in[125]; 
    assign layer_0[3356] = in[680] ^ in[681]; 
    assign layer_0[3357] = ~(in[663] ^ in[501]); 
    assign layer_0[3358] = ~(in[624] | in[606]); 
    assign layer_0[3359] = in[697] & in[710]; 
    assign layer_0[3360] = ~(in[635] ^ in[350]); 
    assign layer_0[3361] = ~(in[731] ^ in[595]); 
    assign layer_0[3362] = in[548] | in[760]; 
    assign layer_0[3363] = ~in[409]; 
    assign layer_0[3364] = in[618] | in[617]; 
    assign layer_0[3365] = in[44] & ~in[298]; 
    assign layer_0[3366] = in[468] & ~in[610]; 
    assign layer_0[3367] = ~(in[634] & in[73]); 
    assign layer_0[3368] = ~in[616] | (in[368] & in[616]); 
    assign layer_0[3369] = ~in[533] | (in[533] & in[553]); 
    assign layer_0[3370] = ~in[488] | (in[488] & in[78]); 
    assign layer_0[3371] = in[148] ^ in[331]; 
    assign layer_0[3372] = ~(in[622] | in[480]); 
    assign layer_0[3373] = in[585] & ~in[284]; 
    assign layer_0[3374] = in[749] | in[582]; 
    assign layer_0[3375] = ~in[88]; 
    assign layer_0[3376] = ~in[252]; 
    assign layer_0[3377] = in[539] ^ in[518]; 
    assign layer_0[3378] = in[536] & in[442]; 
    assign layer_0[3379] = ~(in[682] ^ in[333]); 
    assign layer_0[3380] = in[730] & ~in[620]; 
    assign layer_0[3381] = in[92] & ~in[204]; 
    assign layer_0[3382] = ~(in[338] | in[594]); 
    assign layer_0[3383] = ~(in[282] | in[628]); 
    assign layer_0[3384] = in[435]; 
    assign layer_0[3385] = in[413] ^ in[276]; 
    assign layer_0[3386] = ~(in[259] | in[205]); 
    assign layer_0[3387] = ~(in[649] & in[456]); 
    assign layer_0[3388] = in[87] ^ in[268]; 
    assign layer_0[3389] = ~(in[79] ^ in[709]); 
    assign layer_0[3390] = ~(in[231] & in[573]); 
    assign layer_0[3391] = in[569] & ~in[132]; 
    assign layer_0[3392] = in[45] | in[7]; 
    assign layer_0[3393] = in[34] | in[13]; 
    assign layer_0[3394] = ~(in[460] & in[264]); 
    assign layer_0[3395] = ~(in[651] ^ in[62]); 
    assign layer_0[3396] = ~(in[660] ^ in[161]); 
    assign layer_0[3397] = in[260] ^ in[501]; 
    assign layer_0[3398] = ~(in[754] | in[555]); 
    assign layer_0[3399] = in[343] & in[182]; 
    assign layer_0[3400] = ~(in[414] ^ in[268]); 
    assign layer_0[3401] = in[284] ^ in[364]; 
    assign layer_0[3402] = in[455] ^ in[79]; 
    assign layer_0[3403] = ~(in[412] & in[327]); 
    assign layer_0[3404] = ~(in[563] ^ in[111]); 
    assign layer_0[3405] = in[316] | in[508]; 
    assign layer_0[3406] = ~in[684]; 
    assign layer_0[3407] = ~(in[564] ^ in[683]); 
    assign layer_0[3408] = ~(in[550] ^ in[727]); 
    assign layer_0[3409] = ~in[155] | (in[316] & in[155]); 
    assign layer_0[3410] = in[630] ^ in[201]; 
    assign layer_0[3411] = ~in[380] | (in[5] & in[380]); 
    assign layer_0[3412] = in[350] ^ in[467]; 
    assign layer_0[3413] = 1'b0; 
    assign layer_0[3414] = ~in[637]; 
    assign layer_0[3415] = in[505] ^ in[248]; 
    assign layer_0[3416] = in[652] & ~in[712]; 
    assign layer_0[3417] = ~in[759]; 
    assign layer_0[3418] = ~in[214] | (in[214] & in[661]); 
    assign layer_0[3419] = in[633] ^ in[602]; 
    assign layer_0[3420] = ~in[325]; 
    assign layer_0[3421] = in[319] & in[433]; 
    assign layer_0[3422] = in[60] ^ in[44]; 
    assign layer_0[3423] = in[131] ^ in[742]; 
    assign layer_0[3424] = ~in[375] | (in[475] & in[375]); 
    assign layer_0[3425] = ~in[370] | (in[425] & in[370]); 
    assign layer_0[3426] = in[603]; 
    assign layer_0[3427] = in[250] | in[636]; 
    assign layer_0[3428] = in[573] ^ in[709]; 
    assign layer_0[3429] = ~(in[645] ^ in[275]); 
    assign layer_0[3430] = ~(in[562] | in[34]); 
    assign layer_0[3431] = ~(in[726] ^ in[499]); 
    assign layer_0[3432] = in[246]; 
    assign layer_0[3433] = in[29] | in[650]; 
    assign layer_0[3434] = in[465] ^ in[237]; 
    assign layer_0[3435] = in[692] ^ in[623]; 
    assign layer_0[3436] = in[598] & ~in[665]; 
    assign layer_0[3437] = in[119] & in[267]; 
    assign layer_0[3438] = in[403]; 
    assign layer_0[3439] = in[330] | in[330]; 
    assign layer_0[3440] = in[326]; 
    assign layer_0[3441] = ~(in[508] & in[675]); 
    assign layer_0[3442] = in[311] & ~in[729]; 
    assign layer_0[3443] = in[550] | in[268]; 
    assign layer_0[3444] = ~(in[758] | in[593]); 
    assign layer_0[3445] = ~(in[462] | in[461]); 
    assign layer_0[3446] = ~in[284]; 
    assign layer_0[3447] = in[193] ^ in[418]; 
    assign layer_0[3448] = ~in[598] | (in[307] & in[598]); 
    assign layer_0[3449] = ~(in[613] & in[603]); 
    assign layer_0[3450] = ~in[129]; 
    assign layer_0[3451] = in[655] ^ in[605]; 
    assign layer_0[3452] = in[712] ^ in[360]; 
    assign layer_0[3453] = ~(in[692] ^ in[713]); 
    assign layer_0[3454] = ~(in[596] | in[517]); 
    assign layer_0[3455] = ~(in[518] | in[347]); 
    assign layer_0[3456] = ~(in[77] ^ in[412]); 
    assign layer_0[3457] = ~in[662] | (in[211] & in[662]); 
    assign layer_0[3458] = in[450] & ~in[113]; 
    assign layer_0[3459] = ~(in[84] | in[589]); 
    assign layer_0[3460] = ~in[4] | (in[4] & in[483]); 
    assign layer_0[3461] = ~in[445] | (in[445] & in[178]); 
    assign layer_0[3462] = ~(in[615] ^ in[698]); 
    assign layer_0[3463] = in[230] & ~in[749]; 
    assign layer_0[3464] = ~in[384]; 
    assign layer_0[3465] = ~in[332] | (in[691] & in[332]); 
    assign layer_0[3466] = in[747] ^ in[506]; 
    assign layer_0[3467] = ~(in[607] ^ in[621]); 
    assign layer_0[3468] = ~(in[682] | in[247]); 
    assign layer_0[3469] = in[435] & ~in[536]; 
    assign layer_0[3470] = in[313] ^ in[387]; 
    assign layer_0[3471] = in[473] | in[628]; 
    assign layer_0[3472] = ~in[647] | (in[647] & in[488]); 
    assign layer_0[3473] = 1'b1; 
    assign layer_0[3474] = ~(in[680] & in[616]); 
    assign layer_0[3475] = ~in[325]; 
    assign layer_0[3476] = in[261]; 
    assign layer_0[3477] = in[378] ^ in[694]; 
    assign layer_0[3478] = in[684] & ~in[716]; 
    assign layer_0[3479] = in[710] & ~in[745]; 
    assign layer_0[3480] = in[580] ^ in[142]; 
    assign layer_0[3481] = in[349] ^ in[108]; 
    assign layer_0[3482] = in[696] | in[670]; 
    assign layer_0[3483] = ~in[741]; 
    assign layer_0[3484] = ~(in[602] | in[177]); 
    assign layer_0[3485] = in[762] | in[539]; 
    assign layer_0[3486] = in[68] | in[62]; 
    assign layer_0[3487] = in[592] ^ in[132]; 
    assign layer_0[3488] = in[311] ^ in[35]; 
    assign layer_0[3489] = ~(in[663] ^ in[129]); 
    assign layer_0[3490] = ~(in[210] ^ in[586]); 
    assign layer_0[3491] = ~(in[745] | in[227]); 
    assign layer_0[3492] = in[293] & in[679]; 
    assign layer_0[3493] = ~in[172] | (in[172] & in[320]); 
    assign layer_0[3494] = in[475] ^ in[564]; 
    assign layer_0[3495] = in[347] ^ in[413]; 
    assign layer_0[3496] = in[761] | in[613]; 
    assign layer_0[3497] = in[281] & ~in[761]; 
    assign layer_0[3498] = ~(in[18] ^ in[624]); 
    assign layer_0[3499] = in[28] & ~in[599]; 
    assign layer_0[3500] = in[94] ^ in[358]; 
    assign layer_0[3501] = ~in[392] | (in[392] & in[598]); 
    assign layer_0[3502] = in[417] & ~in[682]; 
    assign layer_0[3503] = ~(in[732] | in[482]); 
    assign layer_0[3504] = ~(in[591] & in[239]); 
    assign layer_0[3505] = ~(in[80] | in[713]); 
    assign layer_0[3506] = in[452] & in[488]; 
    assign layer_0[3507] = in[322] & ~in[363]; 
    assign layer_0[3508] = ~in[309] | (in[646] & in[309]); 
    assign layer_0[3509] = ~in[82] | (in[82] & in[503]); 
    assign layer_0[3510] = in[760] ^ in[611]; 
    assign layer_0[3511] = in[566] | in[483]; 
    assign layer_0[3512] = ~in[579] | (in[579] & in[19]); 
    assign layer_0[3513] = in[628] ^ in[725]; 
    assign layer_0[3514] = ~(in[280] & in[428]); 
    assign layer_0[3515] = in[13] & ~in[710]; 
    assign layer_0[3516] = in[210] | in[3]; 
    assign layer_0[3517] = ~(in[438] ^ in[766]); 
    assign layer_0[3518] = ~in[533] | (in[535] & in[533]); 
    assign layer_0[3519] = ~in[9] | (in[7] & in[9]); 
    assign layer_0[3520] = in[279]; 
    assign layer_0[3521] = in[162] ^ in[599]; 
    assign layer_0[3522] = ~(in[147] | in[690]); 
    assign layer_0[3523] = ~in[421] | (in[668] & in[421]); 
    assign layer_0[3524] = in[656] ^ in[285]; 
    assign layer_0[3525] = in[109] ^ in[688]; 
    assign layer_0[3526] = in[159] & in[243]; 
    assign layer_0[3527] = ~in[665] | (in[41] & in[665]); 
    assign layer_0[3528] = in[277]; 
    assign layer_0[3529] = ~(in[25] & in[760]); 
    assign layer_0[3530] = ~(in[598] | in[551]); 
    assign layer_0[3531] = ~(in[10] ^ in[718]); 
    assign layer_0[3532] = in[458] & in[353]; 
    assign layer_0[3533] = in[564]; 
    assign layer_0[3534] = ~in[134] | (in[134] & in[20]); 
    assign layer_0[3535] = in[342] & ~in[484]; 
    assign layer_0[3536] = ~in[474]; 
    assign layer_0[3537] = ~(in[496] ^ in[420]); 
    assign layer_0[3538] = in[174] ^ in[62]; 
    assign layer_0[3539] = ~(in[760] | in[275]); 
    assign layer_0[3540] = ~(in[502] ^ in[243]); 
    assign layer_0[3541] = in[613] | in[3]; 
    assign layer_0[3542] = ~(in[749] ^ in[760]); 
    assign layer_0[3543] = in[113] | in[624]; 
    assign layer_0[3544] = in[713] & in[709]; 
    assign layer_0[3545] = in[193] | in[746]; 
    assign layer_0[3546] = in[284] ^ in[660]; 
    assign layer_0[3547] = ~in[4] | (in[17] & in[4]); 
    assign layer_0[3548] = ~in[438]; 
    assign layer_0[3549] = ~(in[256] ^ in[153]); 
    assign layer_0[3550] = in[504] & ~in[679]; 
    assign layer_0[3551] = ~(in[623] ^ in[112]); 
    assign layer_0[3552] = in[357]; 
    assign layer_0[3553] = in[173] ^ in[698]; 
    assign layer_0[3554] = in[55] & ~in[674]; 
    assign layer_0[3555] = in[664] ^ in[601]; 
    assign layer_0[3556] = in[572] & in[533]; 
    assign layer_0[3557] = in[358] & ~in[760]; 
    assign layer_0[3558] = ~(in[730] & in[364]); 
    assign layer_0[3559] = in[519] | in[595]; 
    assign layer_0[3560] = ~(in[477] ^ in[724]); 
    assign layer_0[3561] = in[434] ^ in[19]; 
    assign layer_0[3562] = ~in[68]; 
    assign layer_0[3563] = in[121]; 
    assign layer_0[3564] = ~(in[461] ^ in[421]); 
    assign layer_0[3565] = in[404] ^ in[554]; 
    assign layer_0[3566] = in[687] ^ in[647]; 
    assign layer_0[3567] = 1'b1; 
    assign layer_0[3568] = ~(in[759] ^ in[618]); 
    assign layer_0[3569] = in[462] | in[332]; 
    assign layer_0[3570] = in[36] ^ in[699]; 
    assign layer_0[3571] = in[658] ^ in[512]; 
    assign layer_0[3572] = ~in[702] | (in[497] & in[702]); 
    assign layer_0[3573] = ~in[439]; 
    assign layer_0[3574] = ~in[186] | (in[466] & in[186]); 
    assign layer_0[3575] = ~in[493] | (in[493] & in[206]); 
    assign layer_0[3576] = ~(in[291] ^ in[760]); 
    assign layer_0[3577] = ~(in[223] ^ in[266]); 
    assign layer_0[3578] = ~in[498] | (in[372] & in[498]); 
    assign layer_0[3579] = ~(in[499] ^ in[628]); 
    assign layer_0[3580] = in[257] | in[682]; 
    assign layer_0[3581] = ~in[427] | (in[427] & in[46]); 
    assign layer_0[3582] = in[104]; 
    assign layer_0[3583] = ~in[20]; 
    assign layer_0[3584] = ~(in[32] | in[736]); 
    assign layer_0[3585] = ~in[263]; 
    assign layer_0[3586] = ~(in[514] | in[620]); 
    assign layer_0[3587] = ~in[509]; 
    assign layer_0[3588] = ~in[565] | (in[499] & in[565]); 
    assign layer_0[3589] = ~(in[318] ^ in[101]); 
    assign layer_0[3590] = in[281] ^ in[338]; 
    assign layer_0[3591] = in[27] & ~in[658]; 
    assign layer_0[3592] = ~(in[444] ^ in[300]); 
    assign layer_0[3593] = in[18] | in[1]; 
    assign layer_0[3594] = in[340] & ~in[234]; 
    assign layer_0[3595] = ~in[588]; 
    assign layer_0[3596] = ~(in[254] | in[417]); 
    assign layer_0[3597] = ~(in[599] ^ in[198]); 
    assign layer_0[3598] = ~in[441] | (in[723] & in[441]); 
    assign layer_0[3599] = in[436] ^ in[272]; 
    assign layer_0[3600] = ~in[433]; 
    assign layer_0[3601] = in[724]; 
    assign layer_0[3602] = ~(in[486] ^ in[643]); 
    assign layer_0[3603] = in[521] & ~in[434]; 
    assign layer_0[3604] = in[682] & in[645]; 
    assign layer_0[3605] = in[579] & in[440]; 
    assign layer_0[3606] = in[4] & ~in[632]; 
    assign layer_0[3607] = in[263]; 
    assign layer_0[3608] = in[580]; 
    assign layer_0[3609] = ~(in[189] & in[678]); 
    assign layer_0[3610] = in[42] | in[401]; 
    assign layer_0[3611] = ~(in[537] ^ in[697]); 
    assign layer_0[3612] = ~(in[69] ^ in[209]); 
    assign layer_0[3613] = in[535] ^ in[648]; 
    assign layer_0[3614] = in[571] ^ in[523]; 
    assign layer_0[3615] = in[261]; 
    assign layer_0[3616] = ~(in[13] | in[112]); 
    assign layer_0[3617] = in[679] & ~in[158]; 
    assign layer_0[3618] = in[253] & ~in[381]; 
    assign layer_0[3619] = ~(in[45] | in[36]); 
    assign layer_0[3620] = in[709]; 
    assign layer_0[3621] = in[461] | in[365]; 
    assign layer_0[3622] = in[236] ^ in[632]; 
    assign layer_0[3623] = in[760] & ~in[2]; 
    assign layer_0[3624] = ~(in[364] ^ in[698]); 
    assign layer_0[3625] = ~(in[632] ^ in[633]); 
    assign layer_0[3626] = in[168] ^ in[691]; 
    assign layer_0[3627] = ~in[308]; 
    assign layer_0[3628] = ~(in[568] | in[484]); 
    assign layer_0[3629] = ~(in[300] ^ in[512]); 
    assign layer_0[3630] = ~(in[614] ^ in[328]); 
    assign layer_0[3631] = in[253] ^ in[205]; 
    assign layer_0[3632] = in[752] ^ in[309]; 
    assign layer_0[3633] = ~(in[536] ^ in[98]); 
    assign layer_0[3634] = in[696] & in[534]; 
    assign layer_0[3635] = ~in[484] | (in[3] & in[484]); 
    assign layer_0[3636] = ~in[201]; 
    assign layer_0[3637] = ~(in[747] ^ in[8]); 
    assign layer_0[3638] = in[49] | in[466]; 
    assign layer_0[3639] = in[586] ^ in[761]; 
    assign layer_0[3640] = in[397]; 
    assign layer_0[3641] = ~(in[514] | in[490]); 
    assign layer_0[3642] = ~in[680] | (in[680] & in[47]); 
    assign layer_0[3643] = in[323] ^ in[597]; 
    assign layer_0[3644] = in[79] ^ in[23]; 
    assign layer_0[3645] = in[709] ^ in[565]; 
    assign layer_0[3646] = in[755] | in[373]; 
    assign layer_0[3647] = in[252] ^ in[88]; 
    assign layer_0[3648] = ~(in[28] ^ in[296]); 
    assign layer_0[3649] = in[160] & ~in[502]; 
    assign layer_0[3650] = ~in[106] | (in[106] & in[483]); 
    assign layer_0[3651] = ~in[44] | (in[44] & in[745]); 
    assign layer_0[3652] = in[742] & ~in[93]; 
    assign layer_0[3653] = ~(in[355] ^ in[678]); 
    assign layer_0[3654] = in[652]; 
    assign layer_0[3655] = in[355]; 
    assign layer_0[3656] = in[682]; 
    assign layer_0[3657] = ~(in[586] ^ in[597]); 
    assign layer_0[3658] = ~(in[695] ^ in[637]); 
    assign layer_0[3659] = in[712]; 
    assign layer_0[3660] = in[645] ^ in[646]; 
    assign layer_0[3661] = in[454] & ~in[510]; 
    assign layer_0[3662] = ~in[631] | (in[631] & in[570]); 
    assign layer_0[3663] = in[549] & ~in[129]; 
    assign layer_0[3664] = ~(in[568] ^ in[569]); 
    assign layer_0[3665] = ~in[27] | (in[27] & in[353]); 
    assign layer_0[3666] = in[340] | in[498]; 
    assign layer_0[3667] = in[667] ^ in[212]; 
    assign layer_0[3668] = ~(in[159] & in[216]); 
    assign layer_0[3669] = ~in[536]; 
    assign layer_0[3670] = ~in[130] | (in[130] & in[503]); 
    assign layer_0[3671] = ~in[181]; 
    assign layer_0[3672] = ~(in[568] ^ in[745]); 
    assign layer_0[3673] = ~in[103]; 
    assign layer_0[3674] = ~(in[633] ^ in[632]); 
    assign layer_0[3675] = ~(in[757] ^ in[691]); 
    assign layer_0[3676] = ~(in[221] | in[712]); 
    assign layer_0[3677] = in[585] ^ in[564]; 
    assign layer_0[3678] = ~(in[655] | in[75]); 
    assign layer_0[3679] = in[306] | in[10]; 
    assign layer_0[3680] = ~in[681]; 
    assign layer_0[3681] = in[99]; 
    assign layer_0[3682] = ~(in[398] & in[152]); 
    assign layer_0[3683] = in[241] ^ in[2]; 
    assign layer_0[3684] = 1'b0; 
    assign layer_0[3685] = in[584] & ~in[683]; 
    assign layer_0[3686] = in[278] & ~in[710]; 
    assign layer_0[3687] = ~(in[108] | in[576]); 
    assign layer_0[3688] = in[632]; 
    assign layer_0[3689] = ~in[312] | (in[458] & in[312]); 
    assign layer_0[3690] = in[413] ^ in[468]; 
    assign layer_0[3691] = ~in[502]; 
    assign layer_0[3692] = ~in[626] | (in[26] & in[626]); 
    assign layer_0[3693] = in[617]; 
    assign layer_0[3694] = in[388] ^ in[444]; 
    assign layer_0[3695] = in[88] & ~in[718]; 
    assign layer_0[3696] = in[71]; 
    assign layer_0[3697] = in[448]; 
    assign layer_0[3698] = in[66] & in[229]; 
    assign layer_0[3699] = ~in[462] | (in[462] & in[535]); 
    assign layer_0[3700] = in[621] ^ in[500]; 
    assign layer_0[3701] = ~(in[422] | in[193]); 
    assign layer_0[3702] = ~(in[311] & in[167]); 
    assign layer_0[3703] = in[423] & ~in[466]; 
    assign layer_0[3704] = in[332] | in[48]; 
    assign layer_0[3705] = ~(in[503] | in[278]); 
    assign layer_0[3706] = ~(in[264] ^ in[478]); 
    assign layer_0[3707] = in[697] | in[701]; 
    assign layer_0[3708] = ~in[65] | (in[65] & in[671]); 
    assign layer_0[3709] = ~(in[83] ^ in[572]); 
    assign layer_0[3710] = in[519] | in[608]; 
    assign layer_0[3711] = in[615] | in[69]; 
    assign layer_0[3712] = in[391]; 
    assign layer_0[3713] = ~in[340] | (in[340] & in[371]); 
    assign layer_0[3714] = ~in[664]; 
    assign layer_0[3715] = ~(in[441] & in[41]); 
    assign layer_0[3716] = ~(in[262] ^ in[635]); 
    assign layer_0[3717] = in[712] & in[454]; 
    assign layer_0[3718] = ~(in[711] ^ in[365]); 
    assign layer_0[3719] = in[362] | in[547]; 
    assign layer_0[3720] = 1'b1; 
    assign layer_0[3721] = ~(in[90] ^ in[655]); 
    assign layer_0[3722] = ~(in[442] & in[596]); 
    assign layer_0[3723] = in[520] & ~in[554]; 
    assign layer_0[3724] = ~in[698]; 
    assign layer_0[3725] = in[492] | in[492]; 
    assign layer_0[3726] = ~in[549] | (in[549] & in[277]); 
    assign layer_0[3727] = in[603]; 
    assign layer_0[3728] = 1'b0; 
    assign layer_0[3729] = in[617] & ~in[30]; 
    assign layer_0[3730] = in[365]; 
    assign layer_0[3731] = in[201] & ~in[623]; 
    assign layer_0[3732] = in[320] & in[737]; 
    assign layer_0[3733] = in[427]; 
    assign layer_0[3734] = ~in[764]; 
    assign layer_0[3735] = ~in[112] | (in[112] & in[412]); 
    assign layer_0[3736] = in[326] | in[450]; 
    assign layer_0[3737] = in[318] ^ in[356]; 
    assign layer_0[3738] = in[531]; 
    assign layer_0[3739] = 1'b0; 
    assign layer_0[3740] = in[403]; 
    assign layer_0[3741] = ~in[492] | (in[709] & in[492]); 
    assign layer_0[3742] = in[327] ^ in[276]; 
    assign layer_0[3743] = in[63]; 
    assign layer_0[3744] = ~(in[458] | in[61]); 
    assign layer_0[3745] = ~(in[355] ^ in[317]); 
    assign layer_0[3746] = ~in[294]; 
    assign layer_0[3747] = in[468] & ~in[570]; 
    assign layer_0[3748] = 1'b1; 
    assign layer_0[3749] = ~in[279] | (in[279] & in[412]); 
    assign layer_0[3750] = ~in[363] | (in[572] & in[363]); 
    assign layer_0[3751] = in[520]; 
    assign layer_0[3752] = ~(in[758] ^ in[428]); 
    assign layer_0[3753] = ~in[627]; 
    assign layer_0[3754] = ~(in[681] ^ in[569]); 
    assign layer_0[3755] = in[667]; 
    assign layer_0[3756] = ~(in[348] ^ in[615]); 
    assign layer_0[3757] = ~(in[233] ^ in[237]); 
    assign layer_0[3758] = ~in[760] | (in[431] & in[760]); 
    assign layer_0[3759] = ~in[675] | (in[663] & in[675]); 
    assign layer_0[3760] = ~in[552] | (in[552] & in[632]); 
    assign layer_0[3761] = ~in[448]; 
    assign layer_0[3762] = ~(in[143] | in[122]); 
    assign layer_0[3763] = in[474] & in[746]; 
    assign layer_0[3764] = ~in[613] | (in[552] & in[613]); 
    assign layer_0[3765] = ~in[609]; 
    assign layer_0[3766] = in[677] | in[566]; 
    assign layer_0[3767] = ~(in[0] | in[305]); 
    assign layer_0[3768] = ~(in[19] ^ in[503]); 
    assign layer_0[3769] = in[125]; 
    assign layer_0[3770] = in[729] & in[570]; 
    assign layer_0[3771] = ~(in[92] ^ in[682]); 
    assign layer_0[3772] = ~(in[678] ^ in[227]); 
    assign layer_0[3773] = ~(in[326] & in[507]); 
    assign layer_0[3774] = in[460] ^ in[146]; 
    assign layer_0[3775] = ~(in[569] | in[630]); 
    assign layer_0[3776] = in[122]; 
    assign layer_0[3777] = in[293] & in[195]; 
    assign layer_0[3778] = in[663] & ~in[323]; 
    assign layer_0[3779] = ~(in[30] ^ in[192]); 
    assign layer_0[3780] = in[307] & ~in[191]; 
    assign layer_0[3781] = in[706] ^ in[682]; 
    assign layer_0[3782] = ~in[581]; 
    assign layer_0[3783] = ~in[758] | (in[751] & in[758]); 
    assign layer_0[3784] = ~in[635]; 
    assign layer_0[3785] = ~(in[761] ^ in[521]); 
    assign layer_0[3786] = in[440]; 
    assign layer_0[3787] = in[696] & ~in[582]; 
    assign layer_0[3788] = in[710] ^ in[376]; 
    assign layer_0[3789] = ~in[757] | (in[757] & in[366]); 
    assign layer_0[3790] = in[747] & in[357]; 
    assign layer_0[3791] = in[189] & ~in[100]; 
    assign layer_0[3792] = in[710] ^ in[666]; 
    assign layer_0[3793] = in[25] & ~in[35]; 
    assign layer_0[3794] = ~in[679]; 
    assign layer_0[3795] = ~(in[743] ^ in[9]); 
    assign layer_0[3796] = ~(in[555] ^ in[761]); 
    assign layer_0[3797] = ~(in[719] | in[385]); 
    assign layer_0[3798] = ~(in[366] ^ in[81]); 
    assign layer_0[3799] = ~in[308]; 
    assign layer_0[3800] = ~in[586] | (in[586] & in[131]); 
    assign layer_0[3801] = in[57] ^ in[236]; 
    assign layer_0[3802] = ~(in[101] & in[149]); 
    assign layer_0[3803] = in[211] ^ in[81]; 
    assign layer_0[3804] = in[449] & ~in[639]; 
    assign layer_0[3805] = in[381] & in[488]; 
    assign layer_0[3806] = ~in[89] | (in[89] & in[168]); 
    assign layer_0[3807] = ~(in[673] | in[54]); 
    assign layer_0[3808] = in[733]; 
    assign layer_0[3809] = ~(in[158] ^ in[105]); 
    assign layer_0[3810] = ~(in[424] ^ in[452]); 
    assign layer_0[3811] = in[620]; 
    assign layer_0[3812] = ~(in[422] ^ in[81]); 
    assign layer_0[3813] = ~(in[725] ^ in[709]); 
    assign layer_0[3814] = ~(in[459] ^ in[24]); 
    assign layer_0[3815] = ~(in[613] | in[354]); 
    assign layer_0[3816] = in[632] & ~in[471]; 
    assign layer_0[3817] = in[524] & ~in[160]; 
    assign layer_0[3818] = ~(in[326] | in[358]); 
    assign layer_0[3819] = ~in[615]; 
    assign layer_0[3820] = in[4] | in[760]; 
    assign layer_0[3821] = ~in[465] | (in[465] & in[549]); 
    assign layer_0[3822] = ~in[111] | (in[111] & in[600]); 
    assign layer_0[3823] = in[614] & in[500]; 
    assign layer_0[3824] = in[585] ^ in[174]; 
    assign layer_0[3825] = ~in[410] | (in[410] & in[713]); 
    assign layer_0[3826] = in[98] & ~in[488]; 
    assign layer_0[3827] = in[499] & ~in[747]; 
    assign layer_0[3828] = in[56] ^ in[649]; 
    assign layer_0[3829] = ~in[671] | (in[671] & in[127]); 
    assign layer_0[3830] = in[714] | in[646]; 
    assign layer_0[3831] = in[459] ^ in[601]; 
    assign layer_0[3832] = in[93] ^ in[444]; 
    assign layer_0[3833] = ~in[440] | (in[708] & in[440]); 
    assign layer_0[3834] = in[190] | in[418]; 
    assign layer_0[3835] = in[301]; 
    assign layer_0[3836] = in[563] ^ in[713]; 
    assign layer_0[3837] = ~(in[126] ^ in[477]); 
    assign layer_0[3838] = in[743] ^ in[501]; 
    assign layer_0[3839] = ~in[460]; 
    assign layer_0[3840] = ~(in[643] ^ in[571]); 
    assign layer_0[3841] = ~in[653] | (in[653] & in[18]); 
    assign layer_0[3842] = in[622] ^ in[654]; 
    assign layer_0[3843] = ~(in[635] | in[651]); 
    assign layer_0[3844] = ~(in[445] ^ in[703]); 
    assign layer_0[3845] = ~in[501]; 
    assign layer_0[3846] = in[728] ^ in[730]; 
    assign layer_0[3847] = ~(in[597] | in[222]); 
    assign layer_0[3848] = ~in[582]; 
    assign layer_0[3849] = ~in[260] | (in[260] & in[130]); 
    assign layer_0[3850] = ~(in[636] | in[14]); 
    assign layer_0[3851] = ~(in[692] ^ in[605]); 
    assign layer_0[3852] = in[610] & ~in[11]; 
    assign layer_0[3853] = in[583] ^ in[586]; 
    assign layer_0[3854] = in[461] & ~in[550]; 
    assign layer_0[3855] = in[630] | in[146]; 
    assign layer_0[3856] = ~in[68] | (in[68] & in[473]); 
    assign layer_0[3857] = in[677] ^ in[218]; 
    assign layer_0[3858] = in[10] & ~in[396]; 
    assign layer_0[3859] = ~in[373] | (in[757] & in[373]); 
    assign layer_0[3860] = in[710] ^ in[712]; 
    assign layer_0[3861] = ~(in[564] | in[754]); 
    assign layer_0[3862] = in[693] & ~in[499]; 
    assign layer_0[3863] = in[662] & ~in[658]; 
    assign layer_0[3864] = in[480] & ~in[27]; 
    assign layer_0[3865] = ~(in[519] ^ in[436]); 
    assign layer_0[3866] = in[742] & in[88]; 
    assign layer_0[3867] = ~(in[648] ^ in[548]); 
    assign layer_0[3868] = ~(in[600] ^ in[343]); 
    assign layer_0[3869] = in[236] & ~in[434]; 
    assign layer_0[3870] = ~(in[193] ^ in[483]); 
    assign layer_0[3871] = ~(in[367] | in[143]); 
    assign layer_0[3872] = in[214] & ~in[693]; 
    assign layer_0[3873] = ~in[614]; 
    assign layer_0[3874] = ~in[68]; 
    assign layer_0[3875] = ~(in[719] & in[508]); 
    assign layer_0[3876] = ~(in[105] | in[498]); 
    assign layer_0[3877] = in[146]; 
    assign layer_0[3878] = in[441] & ~in[356]; 
    assign layer_0[3879] = ~(in[477] ^ in[280]); 
    assign layer_0[3880] = in[630] ^ in[615]; 
    assign layer_0[3881] = 1'b1; 
    assign layer_0[3882] = in[634] & ~in[762]; 
    assign layer_0[3883] = ~(in[50] & in[321]); 
    assign layer_0[3884] = ~(in[158] & in[381]); 
    assign layer_0[3885] = in[76] ^ in[259]; 
    assign layer_0[3886] = ~(in[658] & in[83]); 
    assign layer_0[3887] = in[154] & in[188]; 
    assign layer_0[3888] = ~(in[8] ^ in[419]); 
    assign layer_0[3889] = ~(in[597] ^ in[164]); 
    assign layer_0[3890] = in[316]; 
    assign layer_0[3891] = ~(in[264] ^ in[262]); 
    assign layer_0[3892] = in[396]; 
    assign layer_0[3893] = ~in[242] | (in[242] & in[501]); 
    assign layer_0[3894] = in[59] | in[620]; 
    assign layer_0[3895] = ~(in[232] ^ in[259]); 
    assign layer_0[3896] = ~(in[646] & in[696]); 
    assign layer_0[3897] = ~(in[738] ^ in[582]); 
    assign layer_0[3898] = in[123] & ~in[320]; 
    assign layer_0[3899] = in[655] ^ in[62]; 
    assign layer_0[3900] = in[549] | in[426]; 
    assign layer_0[3901] = in[203] & ~in[676]; 
    assign layer_0[3902] = ~in[267] | (in[267] & in[590]); 
    assign layer_0[3903] = ~(in[4] ^ in[225]); 
    assign layer_0[3904] = in[366] & ~in[309]; 
    assign layer_0[3905] = ~in[565]; 
    assign layer_0[3906] = in[660] & ~in[410]; 
    assign layer_0[3907] = ~(in[604] ^ in[674]); 
    assign layer_0[3908] = ~(in[622] ^ in[21]); 
    assign layer_0[3909] = ~(in[93] & in[98]); 
    assign layer_0[3910] = ~(in[689] | in[341]); 
    assign layer_0[3911] = in[644] | in[33]; 
    assign layer_0[3912] = 1'b1; 
    assign layer_0[3913] = ~in[342]; 
    assign layer_0[3914] = ~(in[680] ^ in[502]); 
    assign layer_0[3915] = 1'b1; 
    assign layer_0[3916] = in[670] ^ in[631]; 
    assign layer_0[3917] = in[461] & in[242]; 
    assign layer_0[3918] = in[106] ^ in[477]; 
    assign layer_0[3919] = in[712] ^ in[533]; 
    assign layer_0[3920] = ~in[359] | (in[565] & in[359]); 
    assign layer_0[3921] = in[365] | in[89]; 
    assign layer_0[3922] = in[424]; 
    assign layer_0[3923] = in[239] | in[29]; 
    assign layer_0[3924] = in[13] | in[436]; 
    assign layer_0[3925] = 1'b0; 
    assign layer_0[3926] = in[461] ^ in[492]; 
    assign layer_0[3927] = in[381] & in[333]; 
    assign layer_0[3928] = ~(in[332] | in[380]); 
    assign layer_0[3929] = ~(in[491] ^ in[466]); 
    assign layer_0[3930] = in[759] ^ in[667]; 
    assign layer_0[3931] = in[628] & ~in[427]; 
    assign layer_0[3932] = ~in[654] | (in[654] & in[479]); 
    assign layer_0[3933] = in[466] & in[7]; 
    assign layer_0[3934] = ~(in[283] ^ in[413]); 
    assign layer_0[3935] = ~in[370] | (in[370] & in[224]); 
    assign layer_0[3936] = in[276]; 
    assign layer_0[3937] = in[615]; 
    assign layer_0[3938] = in[335] | in[665]; 
    assign layer_0[3939] = in[401] ^ in[296]; 
    assign layer_0[3940] = ~(in[398] ^ in[435]); 
    assign layer_0[3941] = in[498] ^ in[278]; 
    assign layer_0[3942] = in[620] ^ in[358]; 
    assign layer_0[3943] = ~(in[5] ^ in[333]); 
    assign layer_0[3944] = in[574] | in[714]; 
    assign layer_0[3945] = in[611] & ~in[690]; 
    assign layer_0[3946] = in[348] ^ in[662]; 
    assign layer_0[3947] = in[427] ^ in[456]; 
    assign layer_0[3948] = in[730] ^ in[643]; 
    assign layer_0[3949] = ~(in[606] ^ in[241]); 
    assign layer_0[3950] = in[261]; 
    assign layer_0[3951] = in[536] & in[533]; 
    assign layer_0[3952] = in[548] ^ in[298]; 
    assign layer_0[3953] = in[283] & in[429]; 
    assign layer_0[3954] = ~in[152] | (in[187] & in[152]); 
    assign layer_0[3955] = ~in[98] | (in[699] & in[98]); 
    assign layer_0[3956] = in[457] ^ in[706]; 
    assign layer_0[3957] = in[326] ^ in[275]; 
    assign layer_0[3958] = ~in[164] | (in[164] & in[268]); 
    assign layer_0[3959] = ~in[193]; 
    assign layer_0[3960] = ~in[113] | (in[526] & in[113]); 
    assign layer_0[3961] = ~in[54] | (in[64] & in[54]); 
    assign layer_0[3962] = ~in[408]; 
    assign layer_0[3963] = ~(in[428] ^ in[229]); 
    assign layer_0[3964] = in[382] ^ in[223]; 
    assign layer_0[3965] = ~(in[233] ^ in[236]); 
    assign layer_0[3966] = ~in[504] | (in[223] & in[504]); 
    assign layer_0[3967] = 1'b0; 
    assign layer_0[3968] = ~in[669] | (in[669] & in[265]); 
    assign layer_0[3969] = in[292] ^ in[61]; 
    assign layer_0[3970] = in[503]; 
    assign layer_0[3971] = in[44] & ~in[584]; 
    assign layer_0[3972] = ~(in[289] ^ in[397]); 
    assign layer_0[3973] = ~(in[372] ^ in[375]); 
    assign layer_0[3974] = in[463] ^ in[368]; 
    assign layer_0[3975] = ~(in[718] | in[590]); 
    assign layer_0[3976] = ~in[31]; 
    assign layer_0[3977] = ~in[643]; 
    assign layer_0[3978] = in[712] | in[680]; 
    assign layer_0[3979] = in[313] ^ in[331]; 
    assign layer_0[3980] = in[635]; 
    assign layer_0[3981] = in[681] ^ in[246]; 
    assign layer_0[3982] = in[568]; 
    assign layer_0[3983] = ~(in[616] ^ in[569]); 
    assign layer_0[3984] = ~(in[521] ^ in[615]); 
    assign layer_0[3985] = in[312] ^ in[12]; 
    assign layer_0[3986] = in[98] & in[315]; 
    assign layer_0[3987] = ~(in[687] | in[349]); 
    assign layer_0[3988] = in[275] ^ in[461]; 
    assign layer_0[3989] = in[742] ^ in[97]; 
    assign layer_0[3990] = ~in[490]; 
    assign layer_0[3991] = ~(in[586] ^ in[205]); 
    assign layer_0[3992] = ~in[511]; 
    assign layer_0[3993] = in[633] & in[358]; 
    assign layer_0[3994] = in[279] | in[597]; 
    assign layer_0[3995] = ~(in[630] & in[696]); 
    assign layer_0[3996] = in[28] | in[67]; 
    assign layer_0[3997] = in[189] ^ in[553]; 
    assign layer_0[3998] = in[59] & ~in[36]; 
    assign layer_0[3999] = ~(in[574] | in[600]); 
    assign layer_0[4000] = ~(in[713] | in[400]); 
    assign layer_0[4001] = in[401] | in[266]; 
    assign layer_0[4002] = in[362] & in[425]; 
    assign layer_0[4003] = ~in[266] | (in[648] & in[266]); 
    assign layer_0[4004] = ~in[331] | (in[253] & in[331]); 
    assign layer_0[4005] = in[435] & in[654]; 
    assign layer_0[4006] = ~in[165] | (in[165] & in[631]); 
    assign layer_0[4007] = ~(in[549] ^ in[221]); 
    assign layer_0[4008] = ~in[129]; 
    assign layer_0[4009] = ~(in[467] ^ in[482]); 
    assign layer_0[4010] = in[688] ^ in[556]; 
    assign layer_0[4011] = in[527] & ~in[388]; 
    assign layer_0[4012] = ~in[360] | (in[472] & in[360]); 
    assign layer_0[4013] = in[102]; 
    assign layer_0[4014] = in[141] ^ in[428]; 
    assign layer_0[4015] = in[415] ^ in[75]; 
    assign layer_0[4016] = ~(in[298] & in[725]); 
    assign layer_0[4017] = ~(in[66] | in[762]); 
    assign layer_0[4018] = in[267] & in[505]; 
    assign layer_0[4019] = in[42] & in[501]; 
    assign layer_0[4020] = ~in[43] | (in[373] & in[43]); 
    assign layer_0[4021] = ~(in[404] ^ in[242]); 
    assign layer_0[4022] = ~(in[617] ^ in[253]); 
    assign layer_0[4023] = ~(in[284] & in[261]); 
    assign layer_0[4024] = ~(in[209] ^ in[520]); 
    assign layer_0[4025] = 1'b0; 
    assign layer_0[4026] = ~in[574]; 
    assign layer_0[4027] = in[452] ^ in[8]; 
    assign layer_0[4028] = in[583] ^ in[279]; 
    assign layer_0[4029] = ~(in[653] ^ in[337]); 
    assign layer_0[4030] = ~(in[505] ^ in[440]); 
    assign layer_0[4031] = ~in[570] | (in[697] & in[570]); 
    assign layer_0[4032] = ~(in[614] ^ in[692]); 
    assign layer_0[4033] = ~in[591] | (in[591] & in[472]); 
    assign layer_0[4034] = in[34] & ~in[322]; 
    assign layer_0[4035] = ~in[38] | (in[284] & in[38]); 
    assign layer_0[4036] = ~(in[403] ^ in[550]); 
    assign layer_0[4037] = in[548] ^ in[725]; 
    assign layer_0[4038] = in[603] & ~in[694]; 
    assign layer_0[4039] = ~(in[650] | in[651]); 
    assign layer_0[4040] = in[49] ^ in[420]; 
    assign layer_0[4041] = in[12] | in[648]; 
    assign layer_0[4042] = ~(in[693] & in[615]); 
    assign layer_0[4043] = in[358] | in[250]; 
    assign layer_0[4044] = in[647] ^ in[673]; 
    assign layer_0[4045] = ~(in[711] ^ in[324]); 
    assign layer_0[4046] = ~in[395]; 
    assign layer_0[4047] = in[369]; 
    assign layer_0[4048] = ~in[514] | (in[583] & in[514]); 
    assign layer_0[4049] = ~(in[437] & in[508]); 
    assign layer_0[4050] = ~(in[500] & in[19]); 
    assign layer_0[4051] = ~(in[39] & in[421]); 
    assign layer_0[4052] = ~(in[605] ^ in[214]); 
    assign layer_0[4053] = in[91] & in[29]; 
    assign layer_0[4054] = in[195] & ~in[748]; 
    assign layer_0[4055] = ~in[267]; 
    assign layer_0[4056] = ~(in[35] ^ in[207]); 
    assign layer_0[4057] = ~in[154] | (in[154] & in[550]); 
    assign layer_0[4058] = ~in[749] | (in[49] & in[749]); 
    assign layer_0[4059] = in[18]; 
    assign layer_0[4060] = ~(in[350] & in[127]); 
    assign layer_0[4061] = in[189] ^ in[551]; 
    assign layer_0[4062] = ~(in[687] | in[500]); 
    assign layer_0[4063] = ~(in[214] & in[417]); 
    assign layer_0[4064] = ~(in[170] & in[701]); 
    assign layer_0[4065] = ~in[434] | (in[434] & in[349]); 
    assign layer_0[4066] = ~in[490] | (in[174] & in[490]); 
    assign layer_0[4067] = in[685] & ~in[482]; 
    assign layer_0[4068] = ~(in[35] ^ in[275]); 
    assign layer_0[4069] = in[26] & ~in[320]; 
    assign layer_0[4070] = in[81] & in[144]; 
    assign layer_0[4071] = in[758] & ~in[80]; 
    assign layer_0[4072] = ~(in[195] & in[470]); 
    assign layer_0[4073] = in[746] ^ in[615]; 
    assign layer_0[4074] = ~in[344] | (in[344] & in[656]); 
    assign layer_0[4075] = in[248] & ~in[109]; 
    assign layer_0[4076] = 1'b1; 
    assign layer_0[4077] = in[188]; 
    assign layer_0[4078] = ~(in[626] | in[540]); 
    assign layer_0[4079] = in[637] ^ in[718]; 
    assign layer_0[4080] = in[138] & ~in[612]; 
    assign layer_0[4081] = ~(in[74] ^ in[667]); 
    assign layer_0[4082] = ~in[13]; 
    assign layer_0[4083] = in[697] | in[699]; 
    assign layer_0[4084] = ~(in[672] ^ in[203]); 
    assign layer_0[4085] = in[283]; 
    assign layer_0[4086] = ~(in[50] ^ in[695]); 
    assign layer_0[4087] = ~(in[492] ^ in[629]); 
    assign layer_0[4088] = ~(in[466] ^ in[10]); 
    assign layer_0[4089] = ~(in[268] ^ in[82]); 
    assign layer_0[4090] = ~in[95] | (in[95] & in[738]); 
    assign layer_0[4091] = in[731] | in[632]; 
    assign layer_0[4092] = in[76] | in[641]; 
    assign layer_0[4093] = ~(in[533] ^ in[535]); 
    assign layer_0[4094] = ~in[186] | (in[374] & in[186]); 
    assign layer_0[4095] = ~in[291]; 
    assign layer_0[4096] = in[34]; 
    assign layer_0[4097] = in[12]; 
    assign layer_0[4098] = ~in[251]; 
    assign layer_0[4099] = ~in[612] | (in[741] & in[612]); 
    assign layer_0[4100] = in[437] ^ in[298]; 
    assign layer_0[4101] = ~(in[350] & in[634]); 
    assign layer_0[4102] = in[436] ^ in[722]; 
    assign layer_0[4103] = ~in[23]; 
    assign layer_0[4104] = ~(in[267] | in[46]); 
    assign layer_0[4105] = ~in[559]; 
    assign layer_0[4106] = ~(in[318] & in[319]); 
    assign layer_0[4107] = ~in[389] | (in[389] & in[339]); 
    assign layer_0[4108] = ~in[206]; 
    assign layer_0[4109] = ~in[196] | (in[19] & in[196]); 
    assign layer_0[4110] = in[253] ^ in[490]; 
    assign layer_0[4111] = in[749] | in[81]; 
    assign layer_0[4112] = in[58] & in[217]; 
    assign layer_0[4113] = ~in[597] | (in[444] & in[597]); 
    assign layer_0[4114] = ~in[177]; 
    assign layer_0[4115] = in[568] | in[125]; 
    assign layer_0[4116] = ~(in[620] ^ in[276]); 
    assign layer_0[4117] = ~(in[179] & in[82]); 
    assign layer_0[4118] = in[644] ^ in[570]; 
    assign layer_0[4119] = ~(in[682] & in[604]); 
    assign layer_0[4120] = 1'b1; 
    assign layer_0[4121] = in[649]; 
    assign layer_0[4122] = ~(in[282] & in[474]); 
    assign layer_0[4123] = in[292]; 
    assign layer_0[4124] = ~(in[393] | in[112]); 
    assign layer_0[4125] = 1'b0; 
    assign layer_0[4126] = in[156]; 
    assign layer_0[4127] = in[363] ^ in[470]; 
    assign layer_0[4128] = in[538] | in[507]; 
    assign layer_0[4129] = ~(in[555] | in[533]); 
    assign layer_0[4130] = ~(in[579] ^ in[620]); 
    assign layer_0[4131] = ~(in[275] ^ in[659]); 
    assign layer_0[4132] = in[492] | in[687]; 
    assign layer_0[4133] = in[698] & in[403]; 
    assign layer_0[4134] = ~(in[275] | in[722]); 
    assign layer_0[4135] = ~in[244] | (in[244] & in[685]); 
    assign layer_0[4136] = ~(in[666] | in[182]); 
    assign layer_0[4137] = ~(in[696] | in[683]); 
    assign layer_0[4138] = in[283]; 
    assign layer_0[4139] = in[729] & ~in[51]; 
    assign layer_0[4140] = ~in[264] | (in[507] & in[264]); 
    assign layer_0[4141] = ~(in[620] | in[155]); 
    assign layer_0[4142] = in[487]; 
    assign layer_0[4143] = ~(in[616] | in[501]); 
    assign layer_0[4144] = ~(in[749] | in[16]); 
    assign layer_0[4145] = in[742]; 
    assign layer_0[4146] = in[331] | in[725]; 
    assign layer_0[4147] = in[209] & ~in[4]; 
    assign layer_0[4148] = ~in[205] | (in[205] & in[674]); 
    assign layer_0[4149] = in[713] & in[747]; 
    assign layer_0[4150] = ~in[161] | (in[112] & in[161]); 
    assign layer_0[4151] = in[52]; 
    assign layer_0[4152] = ~(in[705] ^ in[688]); 
    assign layer_0[4153] = ~(in[323] & in[120]); 
    assign layer_0[4154] = ~in[50] | (in[623] & in[50]); 
    assign layer_0[4155] = ~(in[62] | in[586]); 
    assign layer_0[4156] = in[537] ^ in[659]; 
    assign layer_0[4157] = ~in[555]; 
    assign layer_0[4158] = ~(in[364] ^ in[332]); 
    assign layer_0[4159] = in[280] & in[691]; 
    assign layer_0[4160] = in[325] | in[643]; 
    assign layer_0[4161] = ~in[283]; 
    assign layer_0[4162] = ~(in[689] | in[261]); 
    assign layer_0[4163] = in[597]; 
    assign layer_0[4164] = in[477] ^ in[468]; 
    assign layer_0[4165] = in[155] & ~in[357]; 
    assign layer_0[4166] = in[354] ^ in[91]; 
    assign layer_0[4167] = in[568]; 
    assign layer_0[4168] = 1'b1; 
    assign layer_0[4169] = in[581] ^ in[262]; 
    assign layer_0[4170] = ~(in[600] | in[499]); 
    assign layer_0[4171] = ~(in[745] ^ in[141]); 
    assign layer_0[4172] = ~(in[536] ^ in[651]); 
    assign layer_0[4173] = ~(in[678] ^ in[690]); 
    assign layer_0[4174] = ~(in[338] | in[759]); 
    assign layer_0[4175] = ~(in[85] | in[389]); 
    assign layer_0[4176] = in[262] & ~in[449]; 
    assign layer_0[4177] = ~(in[348] ^ in[569]); 
    assign layer_0[4178] = in[538] & ~in[179]; 
    assign layer_0[4179] = in[633] ^ in[49]; 
    assign layer_0[4180] = ~(in[293] ^ in[284]); 
    assign layer_0[4181] = in[318]; 
    assign layer_0[4182] = 1'b0; 
    assign layer_0[4183] = ~in[204] | (in[644] & in[204]); 
    assign layer_0[4184] = ~in[345] | (in[4] & in[345]); 
    assign layer_0[4185] = in[23] & ~in[334]; 
    assign layer_0[4186] = ~in[746] | (in[646] & in[746]); 
    assign layer_0[4187] = ~in[355]; 
    assign layer_0[4188] = ~in[365]; 
    assign layer_0[4189] = in[484] ^ in[175]; 
    assign layer_0[4190] = ~in[38] | (in[449] & in[38]); 
    assign layer_0[4191] = in[553] & ~in[481]; 
    assign layer_0[4192] = in[632] ^ in[630]; 
    assign layer_0[4193] = in[388] & ~in[390]; 
    assign layer_0[4194] = ~in[16]; 
    assign layer_0[4195] = ~in[563] | (in[563] & in[176]); 
    assign layer_0[4196] = ~(in[250] ^ in[458]); 
    assign layer_0[4197] = in[0]; 
    assign layer_0[4198] = in[457] ^ in[276]; 
    assign layer_0[4199] = in[664] | in[12]; 
    assign layer_0[4200] = 1'b1; 
    assign layer_0[4201] = ~(in[327] ^ in[19]); 
    assign layer_0[4202] = in[575] & ~in[59]; 
    assign layer_0[4203] = ~(in[644] ^ in[317]); 
    assign layer_0[4204] = in[315] ^ in[505]; 
    assign layer_0[4205] = ~in[427] | (in[724] & in[427]); 
    assign layer_0[4206] = ~(in[237] ^ in[193]); 
    assign layer_0[4207] = in[326] & in[468]; 
    assign layer_0[4208] = in[331] | in[603]; 
    assign layer_0[4209] = ~(in[730] | in[646]); 
    assign layer_0[4210] = ~(in[464] | in[481]); 
    assign layer_0[4211] = 1'b1; 
    assign layer_0[4212] = ~(in[237] & in[598]); 
    assign layer_0[4213] = in[365] | in[95]; 
    assign layer_0[4214] = in[258]; 
    assign layer_0[4215] = in[82] & in[344]; 
    assign layer_0[4216] = in[627] & ~in[282]; 
    assign layer_0[4217] = ~(in[760] & in[427]); 
    assign layer_0[4218] = in[684] & ~in[570]; 
    assign layer_0[4219] = in[741] | in[494]; 
    assign layer_0[4220] = in[260]; 
    assign layer_0[4221] = ~in[273]; 
    assign layer_0[4222] = ~(in[75] ^ in[607]); 
    assign layer_0[4223] = in[535] ^ in[475]; 
    assign layer_0[4224] = ~(in[407] | in[518]); 
    assign layer_0[4225] = in[597] & ~in[714]; 
    assign layer_0[4226] = ~(in[732] | in[732]); 
    assign layer_0[4227] = in[233] ^ in[482]; 
    assign layer_0[4228] = ~(in[713] ^ in[261]); 
    assign layer_0[4229] = ~in[362]; 
    assign layer_0[4230] = in[509] | in[568]; 
    assign layer_0[4231] = ~(in[482] ^ in[609]); 
    assign layer_0[4232] = ~(in[697] ^ in[346]); 
    assign layer_0[4233] = in[98] | in[283]; 
    assign layer_0[4234] = ~in[351] | (in[496] & in[351]); 
    assign layer_0[4235] = ~in[356]; 
    assign layer_0[4236] = ~in[604]; 
    assign layer_0[4237] = in[744] ^ in[745]; 
    assign layer_0[4238] = ~(in[253] | in[680]); 
    assign layer_0[4239] = ~(in[533] ^ in[634]); 
    assign layer_0[4240] = in[141] ^ in[393]; 
    assign layer_0[4241] = in[191] ^ in[604]; 
    assign layer_0[4242] = ~(in[5] & in[141]); 
    assign layer_0[4243] = ~in[210]; 
    assign layer_0[4244] = in[255] ^ in[480]; 
    assign layer_0[4245] = in[670] & ~in[225]; 
    assign layer_0[4246] = ~in[646] | (in[646] & in[605]); 
    assign layer_0[4247] = in[524] | in[260]; 
    assign layer_0[4248] = ~(in[161] ^ in[81]); 
    assign layer_0[4249] = ~(in[488] & in[581]); 
    assign layer_0[4250] = in[92]; 
    assign layer_0[4251] = in[727] ^ in[679]; 
    assign layer_0[4252] = in[118] & ~in[605]; 
    assign layer_0[4253] = ~(in[412] | in[347]); 
    assign layer_0[4254] = in[35] | in[761]; 
    assign layer_0[4255] = ~(in[83] | in[14]); 
    assign layer_0[4256] = in[268] & in[658]; 
    assign layer_0[4257] = ~(in[123] ^ in[459]); 
    assign layer_0[4258] = ~(in[621] | in[316]); 
    assign layer_0[4259] = in[100] ^ in[679]; 
    assign layer_0[4260] = in[619] & ~in[299]; 
    assign layer_0[4261] = in[281] ^ in[263]; 
    assign layer_0[4262] = in[535] | in[587]; 
    assign layer_0[4263] = ~(in[339] ^ in[260]); 
    assign layer_0[4264] = ~in[716] | (in[566] & in[716]); 
    assign layer_0[4265] = in[12] ^ in[742]; 
    assign layer_0[4266] = in[403]; 
    assign layer_0[4267] = ~(in[513] | in[407]); 
    assign layer_0[4268] = ~(in[693] ^ in[344]); 
    assign layer_0[4269] = in[74] & ~in[522]; 
    assign layer_0[4270] = ~(in[249] ^ in[240]); 
    assign layer_0[4271] = in[399] & ~in[31]; 
    assign layer_0[4272] = in[287]; 
    assign layer_0[4273] = in[533] | in[357]; 
    assign layer_0[4274] = in[124]; 
    assign layer_0[4275] = ~(in[335] ^ in[467]); 
    assign layer_0[4276] = in[667] & ~in[549]; 
    assign layer_0[4277] = ~(in[443] ^ in[684]); 
    assign layer_0[4278] = in[761]; 
    assign layer_0[4279] = ~(in[500] & in[307]); 
    assign layer_0[4280] = in[118] & ~in[494]; 
    assign layer_0[4281] = in[739] ^ in[584]; 
    assign layer_0[4282] = ~(in[251] & in[524]); 
    assign layer_0[4283] = in[89] & in[455]; 
    assign layer_0[4284] = ~(in[492] ^ in[82]); 
    assign layer_0[4285] = ~in[113]; 
    assign layer_0[4286] = in[27] ^ in[62]; 
    assign layer_0[4287] = in[355] | in[308]; 
    assign layer_0[4288] = in[352] | in[245]; 
    assign layer_0[4289] = in[731]; 
    assign layer_0[4290] = ~in[298] | (in[298] & in[518]); 
    assign layer_0[4291] = in[54] & ~in[479]; 
    assign layer_0[4292] = ~in[296] | (in[296] & in[597]); 
    assign layer_0[4293] = ~in[665]; 
    assign layer_0[4294] = in[3] ^ in[577]; 
    assign layer_0[4295] = ~(in[761] ^ in[569]); 
    assign layer_0[4296] = ~(in[655] ^ in[71]); 
    assign layer_0[4297] = in[301]; 
    assign layer_0[4298] = in[488] & ~in[612]; 
    assign layer_0[4299] = ~(in[59] | in[704]); 
    assign layer_0[4300] = ~in[696] | (in[696] & in[723]); 
    assign layer_0[4301] = 1'b0; 
    assign layer_0[4302] = ~(in[206] ^ in[399]); 
    assign layer_0[4303] = ~(in[20] | in[12]); 
    assign layer_0[4304] = ~in[308]; 
    assign layer_0[4305] = in[683] | in[82]; 
    assign layer_0[4306] = in[14]; 
    assign layer_0[4307] = ~in[242]; 
    assign layer_0[4308] = ~(in[139] & in[399]); 
    assign layer_0[4309] = ~(in[286] | in[761]); 
    assign layer_0[4310] = in[61] ^ in[636]; 
    assign layer_0[4311] = in[536] & in[252]; 
    assign layer_0[4312] = 1'b1; 
    assign layer_0[4313] = in[566] ^ in[500]; 
    assign layer_0[4314] = in[395] & ~in[260]; 
    assign layer_0[4315] = in[364] ^ in[664]; 
    assign layer_0[4316] = ~in[678]; 
    assign layer_0[4317] = ~in[490]; 
    assign layer_0[4318] = ~(in[206] ^ in[644]); 
    assign layer_0[4319] = in[359]; 
    assign layer_0[4320] = ~in[299]; 
    assign layer_0[4321] = in[3] ^ in[553]; 
    assign layer_0[4322] = in[431]; 
    assign layer_0[4323] = ~(in[359] ^ in[642]); 
    assign layer_0[4324] = ~in[327] | (in[601] & in[327]); 
    assign layer_0[4325] = ~(in[619] ^ in[58]); 
    assign layer_0[4326] = in[202] & ~in[413]; 
    assign layer_0[4327] = in[314] | in[568]; 
    assign layer_0[4328] = ~(in[84] | in[582]); 
    assign layer_0[4329] = ~(in[500] ^ in[614]); 
    assign layer_0[4330] = ~(in[364] ^ in[312]); 
    assign layer_0[4331] = ~in[601]; 
    assign layer_0[4332] = in[604]; 
    assign layer_0[4333] = ~in[758] | (in[27] & in[758]); 
    assign layer_0[4334] = in[745] ^ in[388]; 
    assign layer_0[4335] = ~(in[5] ^ in[491]); 
    assign layer_0[4336] = in[645] ^ in[39]; 
    assign layer_0[4337] = in[447] ^ in[607]; 
    assign layer_0[4338] = ~in[391] | (in[760] & in[391]); 
    assign layer_0[4339] = in[744] & ~in[448]; 
    assign layer_0[4340] = in[568]; 
    assign layer_0[4341] = ~(in[458] ^ in[505]); 
    assign layer_0[4342] = in[364] & ~in[428]; 
    assign layer_0[4343] = in[21] & ~in[735]; 
    assign layer_0[4344] = in[758] ^ in[277]; 
    assign layer_0[4345] = 1'b0; 
    assign layer_0[4346] = in[9] ^ in[159]; 
    assign layer_0[4347] = in[69]; 
    assign layer_0[4348] = in[110] ^ in[709]; 
    assign layer_0[4349] = ~(in[489] ^ in[706]); 
    assign layer_0[4350] = in[674] & ~in[192]; 
    assign layer_0[4351] = ~in[348]; 
    assign layer_0[4352] = in[100] & ~in[300]; 
    assign layer_0[4353] = ~in[178] | (in[178] & in[309]); 
    assign layer_0[4354] = ~in[501] | (in[501] & in[381]); 
    assign layer_0[4355] = ~(in[696] ^ in[57]); 
    assign layer_0[4356] = in[93] & ~in[457]; 
    assign layer_0[4357] = in[588]; 
    assign layer_0[4358] = 1'b1; 
    assign layer_0[4359] = in[639] ^ in[98]; 
    assign layer_0[4360] = in[81] ^ in[275]; 
    assign layer_0[4361] = ~in[454] | (in[454] & in[363]); 
    assign layer_0[4362] = in[566] & ~in[520]; 
    assign layer_0[4363] = ~(in[467] ^ in[468]); 
    assign layer_0[4364] = ~(in[56] & in[5]); 
    assign layer_0[4365] = ~in[57]; 
    assign layer_0[4366] = in[651] ^ in[727]; 
    assign layer_0[4367] = ~(in[338] ^ in[697]); 
    assign layer_0[4368] = ~(in[727] ^ in[744]); 
    assign layer_0[4369] = in[261] | in[491]; 
    assign layer_0[4370] = ~(in[511] & in[679]); 
    assign layer_0[4371] = ~in[492]; 
    assign layer_0[4372] = 1'b1; 
    assign layer_0[4373] = in[277] ^ in[648]; 
    assign layer_0[4374] = ~in[645] | (in[645] & in[550]); 
    assign layer_0[4375] = in[5] & ~in[130]; 
    assign layer_0[4376] = ~in[571]; 
    assign layer_0[4377] = ~(in[125] ^ in[298]); 
    assign layer_0[4378] = in[46] | in[463]; 
    assign layer_0[4379] = in[50] ^ in[467]; 
    assign layer_0[4380] = ~(in[111] | in[737]); 
    assign layer_0[4381] = in[270] & ~in[343]; 
    assign layer_0[4382] = 1'b1; 
    assign layer_0[4383] = in[36] & ~in[602]; 
    assign layer_0[4384] = in[700] ^ in[652]; 
    assign layer_0[4385] = ~(in[371] & in[596]); 
    assign layer_0[4386] = ~in[379] | (in[379] & in[764]); 
    assign layer_0[4387] = in[399] ^ in[631]; 
    assign layer_0[4388] = ~(in[356] & in[440]); 
    assign layer_0[4389] = in[401] & ~in[675]; 
    assign layer_0[4390] = ~(in[356] & in[103]); 
    assign layer_0[4391] = ~in[436] | (in[436] & in[672]); 
    assign layer_0[4392] = in[488] & ~in[661]; 
    assign layer_0[4393] = in[246]; 
    assign layer_0[4394] = in[419] | in[222]; 
    assign layer_0[4395] = in[697] ^ in[85]; 
    assign layer_0[4396] = in[429]; 
    assign layer_0[4397] = ~(in[728] ^ in[299]); 
    assign layer_0[4398] = ~(in[358] ^ in[655]); 
    assign layer_0[4399] = ~(in[147] ^ in[300]); 
    assign layer_0[4400] = in[564] ^ in[618]; 
    assign layer_0[4401] = 1'b0; 
    assign layer_0[4402] = in[649] ^ in[83]; 
    assign layer_0[4403] = ~(in[715] | in[706]); 
    assign layer_0[4404] = in[603] & ~in[379]; 
    assign layer_0[4405] = ~in[506]; 
    assign layer_0[4406] = in[296] ^ in[619]; 
    assign layer_0[4407] = in[194] ^ in[260]; 
    assign layer_0[4408] = in[439] & in[13]; 
    assign layer_0[4409] = ~in[67] | (in[67] & in[46]); 
    assign layer_0[4410] = in[356] ^ in[164]; 
    assign layer_0[4411] = in[266] & in[743]; 
    assign layer_0[4412] = ~in[229] | (in[229] & in[132]); 
    assign layer_0[4413] = ~(in[391] ^ in[682]); 
    assign layer_0[4414] = ~in[39] | (in[638] & in[39]); 
    assign layer_0[4415] = in[459] | in[613]; 
    assign layer_0[4416] = ~(in[668] ^ in[644]); 
    assign layer_0[4417] = in[270] ^ in[337]; 
    assign layer_0[4418] = ~(in[611] ^ in[152]); 
    assign layer_0[4419] = ~(in[440] ^ in[241]); 
    assign layer_0[4420] = in[581] & ~in[195]; 
    assign layer_0[4421] = ~(in[754] ^ in[700]); 
    assign layer_0[4422] = in[638] & ~in[598]; 
    assign layer_0[4423] = ~in[317] | (in[273] & in[317]); 
    assign layer_0[4424] = in[581] | in[25]; 
    assign layer_0[4425] = in[684] ^ in[675]; 
    assign layer_0[4426] = in[199] & ~in[598]; 
    assign layer_0[4427] = ~(in[695] ^ in[331]); 
    assign layer_0[4428] = in[614] ^ in[296]; 
    assign layer_0[4429] = in[580] ^ in[93]; 
    assign layer_0[4430] = in[34] & ~in[226]; 
    assign layer_0[4431] = in[548]; 
    assign layer_0[4432] = ~in[9] | (in[374] & in[9]); 
    assign layer_0[4433] = in[159] ^ in[176]; 
    assign layer_0[4434] = ~(in[433] ^ in[356]); 
    assign layer_0[4435] = ~(in[189] ^ in[136]); 
    assign layer_0[4436] = ~(in[30] ^ in[40]); 
    assign layer_0[4437] = in[532] & ~in[305]; 
    assign layer_0[4438] = in[53] ^ in[532]; 
    assign layer_0[4439] = in[207]; 
    assign layer_0[4440] = ~(in[27] ^ in[509]); 
    assign layer_0[4441] = in[72] & ~in[52]; 
    assign layer_0[4442] = in[763] ^ in[617]; 
    assign layer_0[4443] = in[500] ^ in[680]; 
    assign layer_0[4444] = ~(in[715] | in[446]); 
    assign layer_0[4445] = ~in[427] | (in[427] & in[582]); 
    assign layer_0[4446] = ~in[410]; 
    assign layer_0[4447] = ~(in[296] ^ in[3]); 
    assign layer_0[4448] = in[83] & in[113]; 
    assign layer_0[4449] = ~(in[364] ^ in[316]); 
    assign layer_0[4450] = ~(in[605] ^ in[649]); 
    assign layer_0[4451] = ~(in[69] | in[55]); 
    assign layer_0[4452] = ~in[98]; 
    assign layer_0[4453] = in[299] & ~in[491]; 
    assign layer_0[4454] = in[51]; 
    assign layer_0[4455] = in[551] & ~in[507]; 
    assign layer_0[4456] = in[78] & ~in[630]; 
    assign layer_0[4457] = ~in[252]; 
    assign layer_0[4458] = in[143] & ~in[368]; 
    assign layer_0[4459] = in[520] ^ in[599]; 
    assign layer_0[4460] = in[292] ^ in[127]; 
    assign layer_0[4461] = ~in[324]; 
    assign layer_0[4462] = ~(in[156] & in[64]); 
    assign layer_0[4463] = ~(in[313] ^ in[312]); 
    assign layer_0[4464] = 1'b1; 
    assign layer_0[4465] = in[299] & ~in[538]; 
    assign layer_0[4466] = in[426] & in[377]; 
    assign layer_0[4467] = ~in[676] | (in[529] & in[676]); 
    assign layer_0[4468] = ~in[52]; 
    assign layer_0[4469] = in[54] & ~in[84]; 
    assign layer_0[4470] = in[610] | in[562]; 
    assign layer_0[4471] = ~in[710] | (in[710] & in[275]); 
    assign layer_0[4472] = ~in[309] | (in[309] & in[614]); 
    assign layer_0[4473] = in[726]; 
    assign layer_0[4474] = ~in[671] | (in[60] & in[671]); 
    assign layer_0[4475] = in[651] & ~in[293]; 
    assign layer_0[4476] = ~in[3] | (in[610] & in[3]); 
    assign layer_0[4477] = in[508] ^ in[349]; 
    assign layer_0[4478] = ~(in[737] ^ in[5]); 
    assign layer_0[4479] = in[63] ^ in[646]; 
    assign layer_0[4480] = in[687] | in[672]; 
    assign layer_0[4481] = ~(in[429] | in[577]); 
    assign layer_0[4482] = in[95] & ~in[590]; 
    assign layer_0[4483] = in[585] ^ in[291]; 
    assign layer_0[4484] = ~in[130]; 
    assign layer_0[4485] = ~(in[442] & in[423]); 
    assign layer_0[4486] = in[201] ^ in[655]; 
    assign layer_0[4487] = ~in[57]; 
    assign layer_0[4488] = ~in[641] | (in[641] & in[319]); 
    assign layer_0[4489] = ~(in[597] ^ in[490]); 
    assign layer_0[4490] = 1'b1; 
    assign layer_0[4491] = ~(in[34] ^ in[397]); 
    assign layer_0[4492] = ~in[405]; 
    assign layer_0[4493] = in[484] ^ in[444]; 
    assign layer_0[4494] = ~in[315]; 
    assign layer_0[4495] = ~(in[730] & in[539]); 
    assign layer_0[4496] = ~in[244] | (in[618] & in[244]); 
    assign layer_0[4497] = in[301] | in[697]; 
    assign layer_0[4498] = in[654]; 
    assign layer_0[4499] = ~in[501] | (in[631] & in[501]); 
    assign layer_0[4500] = in[286] | in[251]; 
    assign layer_0[4501] = in[179] & ~in[681]; 
    assign layer_0[4502] = in[610] ^ in[92]; 
    assign layer_0[4503] = ~(in[332] ^ in[175]); 
    assign layer_0[4504] = 1'b0; 
    assign layer_0[4505] = in[716] ^ in[662]; 
    assign layer_0[4506] = ~in[682] | (in[682] & in[687]); 
    assign layer_0[4507] = in[106] ^ in[275]; 
    assign layer_0[4508] = in[230] & in[764]; 
    assign layer_0[4509] = ~in[447] | (in[319] & in[447]); 
    assign layer_0[4510] = in[161] & ~in[226]; 
    assign layer_0[4511] = in[387] ^ in[451]; 
    assign layer_0[4512] = in[98] | in[275]; 
    assign layer_0[4513] = ~(in[242] & in[618]); 
    assign layer_0[4514] = ~in[322] | (in[322] & in[348]); 
    assign layer_0[4515] = ~(in[432] | in[613]); 
    assign layer_0[4516] = ~(in[534] ^ in[618]); 
    assign layer_0[4517] = in[708] ^ in[628]; 
    assign layer_0[4518] = in[330] & ~in[313]; 
    assign layer_0[4519] = ~in[37]; 
    assign layer_0[4520] = ~(in[467] ^ in[241]); 
    assign layer_0[4521] = ~(in[151] ^ in[730]); 
    assign layer_0[4522] = in[164] & ~in[300]; 
    assign layer_0[4523] = ~(in[282] ^ in[595]); 
    assign layer_0[4524] = ~in[205] | (in[205] & in[51]); 
    assign layer_0[4525] = ~(in[235] ^ in[599]); 
    assign layer_0[4526] = 1'b1; 
    assign layer_0[4527] = in[331]; 
    assign layer_0[4528] = in[526] ^ in[632]; 
    assign layer_0[4529] = in[252] ^ in[264]; 
    assign layer_0[4530] = in[765] ^ in[250]; 
    assign layer_0[4531] = in[355] & in[69]; 
    assign layer_0[4532] = ~(in[210] ^ in[369]); 
    assign layer_0[4533] = ~in[190]; 
    assign layer_0[4534] = in[149] | in[149]; 
    assign layer_0[4535] = in[373]; 
    assign layer_0[4536] = ~in[470] | (in[492] & in[470]); 
    assign layer_0[4537] = in[430] ^ in[122]; 
    assign layer_0[4538] = in[417] & ~in[128]; 
    assign layer_0[4539] = ~(in[2] | in[283]); 
    assign layer_0[4540] = ~in[145]; 
    assign layer_0[4541] = in[603]; 
    assign layer_0[4542] = ~in[326] | (in[542] & in[326]); 
    assign layer_0[4543] = ~(in[412] & in[349]); 
    assign layer_0[4544] = ~(in[637] ^ in[587]); 
    assign layer_0[4545] = in[267] | in[459]; 
    assign layer_0[4546] = in[118] & in[538]; 
    assign layer_0[4547] = in[698] | in[448]; 
    assign layer_0[4548] = in[29] ^ in[404]; 
    assign layer_0[4549] = ~(in[682] | in[585]); 
    assign layer_0[4550] = in[53]; 
    assign layer_0[4551] = ~in[659] | (in[253] & in[659]); 
    assign layer_0[4552] = in[277]; 
    assign layer_0[4553] = ~in[632] | (in[311] & in[632]); 
    assign layer_0[4554] = ~in[633]; 
    assign layer_0[4555] = in[209] | in[113]; 
    assign layer_0[4556] = ~(in[738] ^ in[651]); 
    assign layer_0[4557] = ~(in[385] ^ in[685]); 
    assign layer_0[4558] = ~(in[402] ^ in[263]); 
    assign layer_0[4559] = in[412] ^ in[731]; 
    assign layer_0[4560] = in[651] & ~in[620]; 
    assign layer_0[4561] = ~(in[513] | in[79]); 
    assign layer_0[4562] = in[747] ^ in[92]; 
    assign layer_0[4563] = ~(in[621] ^ in[333]); 
    assign layer_0[4564] = in[444]; 
    assign layer_0[4565] = ~in[376] | (in[376] & in[96]); 
    assign layer_0[4566] = in[666] ^ in[727]; 
    assign layer_0[4567] = ~(in[692] ^ in[518]); 
    assign layer_0[4568] = ~(in[342] | in[6]); 
    assign layer_0[4569] = ~(in[490] ^ in[740]); 
    assign layer_0[4570] = ~(in[351] ^ in[573]); 
    assign layer_0[4571] = in[415] & ~in[550]; 
    assign layer_0[4572] = ~(in[244] & in[435]); 
    assign layer_0[4573] = ~in[61] | (in[61] & in[673]); 
    assign layer_0[4574] = ~(in[645] & in[694]); 
    assign layer_0[4575] = in[758]; 
    assign layer_0[4576] = in[536]; 
    assign layer_0[4577] = ~in[143] | (in[381] & in[143]); 
    assign layer_0[4578] = in[604] ^ in[101]; 
    assign layer_0[4579] = in[613] ^ in[571]; 
    assign layer_0[4580] = ~in[758] | (in[108] & in[758]); 
    assign layer_0[4581] = in[404] ^ in[290]; 
    assign layer_0[4582] = in[660] ^ in[508]; 
    assign layer_0[4583] = in[84] | in[2]; 
    assign layer_0[4584] = in[675] & ~in[744]; 
    assign layer_0[4585] = in[472] & ~in[94]; 
    assign layer_0[4586] = ~(in[65] | in[321]); 
    assign layer_0[4587] = ~in[767]; 
    assign layer_0[4588] = ~in[406] | (in[397] & in[406]); 
    assign layer_0[4589] = in[467] & ~in[348]; 
    assign layer_0[4590] = in[142]; 
    assign layer_0[4591] = ~(in[719] ^ in[733]); 
    assign layer_0[4592] = ~(in[364] & in[43]); 
    assign layer_0[4593] = in[322] | in[477]; 
    assign layer_0[4594] = in[253] | in[663]; 
    assign layer_0[4595] = in[619] & ~in[53]; 
    assign layer_0[4596] = ~in[455] | (in[455] & in[680]); 
    assign layer_0[4597] = in[5] & ~in[594]; 
    assign layer_0[4598] = in[627] & in[138]; 
    assign layer_0[4599] = in[372] & ~in[179]; 
    assign layer_0[4600] = in[3] & ~in[651]; 
    assign layer_0[4601] = ~(in[486] ^ in[27]); 
    assign layer_0[4602] = 1'b1; 
    assign layer_0[4603] = ~(in[291] & in[745]); 
    assign layer_0[4604] = ~in[645] | (in[645] & in[762]); 
    assign layer_0[4605] = in[147] & ~in[657]; 
    assign layer_0[4606] = ~(in[210] & in[323]); 
    assign layer_0[4607] = in[19]; 
    assign layer_0[4608] = ~in[140] | (in[449] & in[140]); 
    assign layer_0[4609] = ~in[220] | (in[220] & in[388]); 
    assign layer_0[4610] = ~in[741] | (in[261] & in[741]); 
    assign layer_0[4611] = ~(in[161] ^ in[378]); 
    assign layer_0[4612] = ~in[519]; 
    assign layer_0[4613] = in[689] & in[628]; 
    assign layer_0[4614] = ~(in[46] ^ in[106]); 
    assign layer_0[4615] = ~in[319] | (in[319] & in[619]); 
    assign layer_0[4616] = in[311]; 
    assign layer_0[4617] = ~in[552] | (in[718] & in[552]); 
    assign layer_0[4618] = in[131] & in[588]; 
    assign layer_0[4619] = in[431] ^ in[303]; 
    assign layer_0[4620] = ~(in[486] | in[599]); 
    assign layer_0[4621] = in[490] ^ in[177]; 
    assign layer_0[4622] = in[40] | in[69]; 
    assign layer_0[4623] = ~in[748]; 
    assign layer_0[4624] = in[436] & ~in[345]; 
    assign layer_0[4625] = in[603] ^ in[583]; 
    assign layer_0[4626] = ~(in[404] | in[593]); 
    assign layer_0[4627] = ~(in[182] & in[651]); 
    assign layer_0[4628] = in[335]; 
    assign layer_0[4629] = ~in[106]; 
    assign layer_0[4630] = ~(in[363] ^ in[171]); 
    assign layer_0[4631] = ~(in[663] ^ in[709]); 
    assign layer_0[4632] = ~(in[411] | in[548]); 
    assign layer_0[4633] = in[649] ^ in[731]; 
    assign layer_0[4634] = in[405] & in[693]; 
    assign layer_0[4635] = in[590] & ~in[370]; 
    assign layer_0[4636] = in[617] ^ in[731]; 
    assign layer_0[4637] = in[756] ^ in[763]; 
    assign layer_0[4638] = ~(in[647] | in[645]); 
    assign layer_0[4639] = in[376] & ~in[338]; 
    assign layer_0[4640] = in[393]; 
    assign layer_0[4641] = ~(in[587] ^ in[67]); 
    assign layer_0[4642] = ~(in[320] | in[762]); 
    assign layer_0[4643] = ~in[473] | (in[763] & in[473]); 
    assign layer_0[4644] = in[428] | in[444]; 
    assign layer_0[4645] = in[36] | in[620]; 
    assign layer_0[4646] = ~in[47] | (in[47] & in[715]); 
    assign layer_0[4647] = in[521] | in[550]; 
    assign layer_0[4648] = ~(in[708] | in[501]); 
    assign layer_0[4649] = ~(in[332] | in[596]); 
    assign layer_0[4650] = ~in[266]; 
    assign layer_0[4651] = ~(in[301] | in[370]); 
    assign layer_0[4652] = in[364]; 
    assign layer_0[4653] = ~(in[316] ^ in[92]); 
    assign layer_0[4654] = in[174] | in[570]; 
    assign layer_0[4655] = in[223] & ~in[70]; 
    assign layer_0[4656] = ~in[398] | (in[37] & in[398]); 
    assign layer_0[4657] = ~in[666] | (in[484] & in[666]); 
    assign layer_0[4658] = in[237] ^ in[372]; 
    assign layer_0[4659] = in[707] ^ in[698]; 
    assign layer_0[4660] = ~(in[604] | in[537]); 
    assign layer_0[4661] = in[340] & ~in[64]; 
    assign layer_0[4662] = ~(in[586] ^ in[86]); 
    assign layer_0[4663] = in[344] ^ in[705]; 
    assign layer_0[4664] = ~(in[570] ^ in[219]); 
    assign layer_0[4665] = in[81] | in[308]; 
    assign layer_0[4666] = in[646] | in[327]; 
    assign layer_0[4667] = ~(in[501] ^ in[388]); 
    assign layer_0[4668] = ~(in[12] ^ in[377]); 
    assign layer_0[4669] = ~in[296] | (in[277] & in[296]); 
    assign layer_0[4670] = in[535] & ~in[220]; 
    assign layer_0[4671] = in[172] ^ in[35]; 
    assign layer_0[4672] = in[522] & ~in[179]; 
    assign layer_0[4673] = ~(in[330] ^ in[625]); 
    assign layer_0[4674] = in[243] & ~in[492]; 
    assign layer_0[4675] = in[546] & in[767]; 
    assign layer_0[4676] = ~(in[106] & in[528]); 
    assign layer_0[4677] = ~(in[568] | in[65]); 
    assign layer_0[4678] = ~in[602]; 
    assign layer_0[4679] = ~in[435] | (in[435] & in[448]); 
    assign layer_0[4680] = ~(in[219] ^ in[681]); 
    assign layer_0[4681] = ~in[207]; 
    assign layer_0[4682] = ~(in[460] ^ in[555]); 
    assign layer_0[4683] = ~(in[248] & in[683]); 
    assign layer_0[4684] = ~in[569] | (in[701] & in[569]); 
    assign layer_0[4685] = in[329] & ~in[517]; 
    assign layer_0[4686] = in[347]; 
    assign layer_0[4687] = ~in[679] | (in[756] & in[679]); 
    assign layer_0[4688] = 1'b0; 
    assign layer_0[4689] = in[760] | in[695]; 
    assign layer_0[4690] = in[59] ^ in[677]; 
    assign layer_0[4691] = in[587] ^ in[373]; 
    assign layer_0[4692] = in[185] ^ in[101]; 
    assign layer_0[4693] = in[95] & ~in[576]; 
    assign layer_0[4694] = in[399] & ~in[98]; 
    assign layer_0[4695] = in[373] ^ in[360]; 
    assign layer_0[4696] = ~(in[584] & in[394]); 
    assign layer_0[4697] = ~(in[195] ^ in[19]); 
    assign layer_0[4698] = ~(in[135] & in[68]); 
    assign layer_0[4699] = in[583] ^ in[210]; 
    assign layer_0[4700] = in[581] ^ in[583]; 
    assign layer_0[4701] = ~in[196] | (in[196] & in[652]); 
    assign layer_0[4702] = in[707] & in[565]; 
    assign layer_0[4703] = ~in[451] | (in[451] & in[521]); 
    assign layer_0[4704] = in[482]; 
    assign layer_0[4705] = in[554] ^ in[115]; 
    assign layer_0[4706] = in[633]; 
    assign layer_0[4707] = in[69]; 
    assign layer_0[4708] = ~in[728] | (in[728] & in[580]); 
    assign layer_0[4709] = ~(in[384] & in[459]); 
    assign layer_0[4710] = ~in[49]; 
    assign layer_0[4711] = in[267]; 
    assign layer_0[4712] = in[549]; 
    assign layer_0[4713] = ~(in[499] & in[93]); 
    assign layer_0[4714] = in[382] ^ in[358]; 
    assign layer_0[4715] = ~(in[70] ^ in[714]); 
    assign layer_0[4716] = in[148] | in[121]; 
    assign layer_0[4717] = in[162] & ~in[652]; 
    assign layer_0[4718] = in[649] ^ in[648]; 
    assign layer_0[4719] = ~(in[254] ^ in[432]); 
    assign layer_0[4720] = in[458] ^ in[71]; 
    assign layer_0[4721] = in[316] & ~in[236]; 
    assign layer_0[4722] = in[84] ^ in[649]; 
    assign layer_0[4723] = in[116] & ~in[721]; 
    assign layer_0[4724] = in[67] | in[721]; 
    assign layer_0[4725] = ~in[601]; 
    assign layer_0[4726] = in[487] & ~in[421]; 
    assign layer_0[4727] = in[251] & ~in[613]; 
    assign layer_0[4728] = ~in[62]; 
    assign layer_0[4729] = in[636]; 
    assign layer_0[4730] = in[225] & ~in[338]; 
    assign layer_0[4731] = ~(in[416] & in[330]); 
    assign layer_0[4732] = ~(in[614] ^ in[71]); 
    assign layer_0[4733] = ~(in[467] ^ in[178]); 
    assign layer_0[4734] = ~in[682] | (in[682] & in[205]); 
    assign layer_0[4735] = ~(in[376] ^ in[699]); 
    assign layer_0[4736] = ~(in[582] ^ in[518]); 
    assign layer_0[4737] = in[503] ^ in[478]; 
    assign layer_0[4738] = in[359] & ~in[166]; 
    assign layer_0[4739] = ~in[525] | (in[525] & in[195]); 
    assign layer_0[4740] = in[178] ^ in[146]; 
    assign layer_0[4741] = in[645] ^ in[439]; 
    assign layer_0[4742] = ~in[503]; 
    assign layer_0[4743] = ~(in[240] | in[368]); 
    assign layer_0[4744] = ~in[431] | (in[26] & in[431]); 
    assign layer_0[4745] = in[663]; 
    assign layer_0[4746] = ~(in[269] ^ in[759]); 
    assign layer_0[4747] = in[453] & ~in[365]; 
    assign layer_0[4748] = ~(in[501] ^ in[548]); 
    assign layer_0[4749] = ~in[335] | (in[335] & in[588]); 
    assign layer_0[4750] = in[618] & ~in[762]; 
    assign layer_0[4751] = ~(in[551] ^ in[460]); 
    assign layer_0[4752] = in[577] ^ in[423]; 
    assign layer_0[4753] = in[132] & in[8]; 
    assign layer_0[4754] = in[656] | in[622]; 
    assign layer_0[4755] = ~in[532] | (in[130] & in[532]); 
    assign layer_0[4756] = ~in[602]; 
    assign layer_0[4757] = ~(in[94] ^ in[284]); 
    assign layer_0[4758] = ~(in[725] ^ in[538]); 
    assign layer_0[4759] = in[115] & in[236]; 
    assign layer_0[4760] = ~(in[677] ^ in[744]); 
    assign layer_0[4761] = in[298] ^ in[355]; 
    assign layer_0[4762] = ~(in[604] ^ in[724]); 
    assign layer_0[4763] = in[34] & ~in[463]; 
    assign layer_0[4764] = in[412] & ~in[127]; 
    assign layer_0[4765] = ~in[555]; 
    assign layer_0[4766] = ~in[101] | (in[306] & in[101]); 
    assign layer_0[4767] = in[343] & ~in[365]; 
    assign layer_0[4768] = ~in[484]; 
    assign layer_0[4769] = ~in[279] | (in[682] & in[279]); 
    assign layer_0[4770] = ~in[212] | (in[112] & in[212]); 
    assign layer_0[4771] = 1'b1; 
    assign layer_0[4772] = in[709]; 
    assign layer_0[4773] = ~(in[307] ^ in[371]); 
    assign layer_0[4774] = in[603] & in[653]; 
    assign layer_0[4775] = ~in[380]; 
    assign layer_0[4776] = in[295] ^ in[650]; 
    assign layer_0[4777] = in[445] ^ in[760]; 
    assign layer_0[4778] = in[584] ^ in[614]; 
    assign layer_0[4779] = ~(in[640] ^ in[520]); 
    assign layer_0[4780] = ~(in[159] ^ in[301]); 
    assign layer_0[4781] = ~in[38] | (in[38] & in[572]); 
    assign layer_0[4782] = in[705] ^ in[755]; 
    assign layer_0[4783] = in[2]; 
    assign layer_0[4784] = ~in[419]; 
    assign layer_0[4785] = ~(in[385] & in[341]); 
    assign layer_0[4786] = ~in[308] | (in[308] & in[306]); 
    assign layer_0[4787] = ~in[714] | (in[188] & in[714]); 
    assign layer_0[4788] = in[655] | in[639]; 
    assign layer_0[4789] = in[283]; 
    assign layer_0[4790] = in[444] & in[50]; 
    assign layer_0[4791] = in[46]; 
    assign layer_0[4792] = ~(in[472] ^ in[685]); 
    assign layer_0[4793] = ~in[26] | (in[331] & in[26]); 
    assign layer_0[4794] = ~(in[674] & in[702]); 
    assign layer_0[4795] = in[295] ^ in[253]; 
    assign layer_0[4796] = in[601]; 
    assign layer_0[4797] = ~in[299] | (in[522] & in[299]); 
    assign layer_0[4798] = ~in[757]; 
    assign layer_0[4799] = in[595] ^ in[723]; 
    assign layer_0[4800] = ~(in[666] | in[492]); 
    assign layer_0[4801] = in[535] & ~in[630]; 
    assign layer_0[4802] = ~in[172] | (in[501] & in[172]); 
    assign layer_0[4803] = in[675] | in[183]; 
    assign layer_0[4804] = 1'b0; 
    assign layer_0[4805] = ~(in[93] ^ in[243]); 
    assign layer_0[4806] = in[694]; 
    assign layer_0[4807] = in[653] & ~in[97]; 
    assign layer_0[4808] = in[125] | in[580]; 
    assign layer_0[4809] = in[570] ^ in[536]; 
    assign layer_0[4810] = in[93] & in[466]; 
    assign layer_0[4811] = ~in[141] | (in[539] & in[141]); 
    assign layer_0[4812] = in[497] | in[629]; 
    assign layer_0[4813] = in[11] ^ in[759]; 
    assign layer_0[4814] = in[758]; 
    assign layer_0[4815] = in[95]; 
    assign layer_0[4816] = in[714] ^ in[281]; 
    assign layer_0[4817] = in[749] ^ in[710]; 
    assign layer_0[4818] = in[242] ^ in[484]; 
    assign layer_0[4819] = in[241] | in[462]; 
    assign layer_0[4820] = ~(in[694] & in[693]); 
    assign layer_0[4821] = ~in[492] | (in[579] & in[492]); 
    assign layer_0[4822] = in[613]; 
    assign layer_0[4823] = in[97] & ~in[326]; 
    assign layer_0[4824] = in[643] ^ in[506]; 
    assign layer_0[4825] = in[574] | in[233]; 
    assign layer_0[4826] = ~(in[179] ^ in[613]); 
    assign layer_0[4827] = in[401] | in[68]; 
    assign layer_0[4828] = in[708] & ~in[704]; 
    assign layer_0[4829] = ~in[646]; 
    assign layer_0[4830] = in[30]; 
    assign layer_0[4831] = ~in[685] | (in[367] & in[685]); 
    assign layer_0[4832] = ~(in[595] | in[347]); 
    assign layer_0[4833] = ~(in[310] ^ in[4]); 
    assign layer_0[4834] = ~in[29] | (in[29] & in[626]); 
    assign layer_0[4835] = in[136]; 
    assign layer_0[4836] = ~(in[98] & in[226]); 
    assign layer_0[4837] = ~(in[615] ^ in[603]); 
    assign layer_0[4838] = in[30]; 
    assign layer_0[4839] = in[62] ^ in[497]; 
    assign layer_0[4840] = in[686]; 
    assign layer_0[4841] = ~(in[636] ^ in[284]); 
    assign layer_0[4842] = 1'b0; 
    assign layer_0[4843] = in[402]; 
    assign layer_0[4844] = ~(in[635] | in[20]); 
    assign layer_0[4845] = ~in[185] | (in[63] & in[185]); 
    assign layer_0[4846] = ~(in[463] & in[673]); 
    assign layer_0[4847] = ~(in[423] & in[595]); 
    assign layer_0[4848] = in[414] & ~in[45]; 
    assign layer_0[4849] = in[245] ^ in[603]; 
    assign layer_0[4850] = ~in[727] | (in[727] & in[404]); 
    assign layer_0[4851] = ~(in[636] & in[3]); 
    assign layer_0[4852] = ~in[67] | (in[275] & in[67]); 
    assign layer_0[4853] = in[483] ^ in[293]; 
    assign layer_0[4854] = in[456] & in[627]; 
    assign layer_0[4855] = ~in[13] | (in[13] & in[405]); 
    assign layer_0[4856] = ~in[297]; 
    assign layer_0[4857] = in[100] & ~in[189]; 
    assign layer_0[4858] = in[5] | in[643]; 
    assign layer_0[4859] = ~(in[537] | in[536]); 
    assign layer_0[4860] = ~in[279]; 
    assign layer_0[4861] = ~in[727]; 
    assign layer_0[4862] = ~(in[744] & in[618]); 
    assign layer_0[4863] = ~(in[267] | in[459]); 
    assign layer_0[4864] = ~in[28] | (in[28] & in[506]); 
    assign layer_0[4865] = in[691]; 
    assign layer_0[4866] = in[460]; 
    assign layer_0[4867] = ~in[9]; 
    assign layer_0[4868] = ~in[341] | (in[683] & in[341]); 
    assign layer_0[4869] = in[469]; 
    assign layer_0[4870] = ~(in[650] ^ in[459]); 
    assign layer_0[4871] = ~(in[446] | in[191]); 
    assign layer_0[4872] = in[567] ^ in[262]; 
    assign layer_0[4873] = ~(in[694] & in[691]); 
    assign layer_0[4874] = ~(in[554] ^ in[533]); 
    assign layer_0[4875] = ~in[408] | (in[173] & in[408]); 
    assign layer_0[4876] = ~in[374] | (in[374] & in[538]); 
    assign layer_0[4877] = in[19] ^ in[264]; 
    assign layer_0[4878] = in[82]; 
    assign layer_0[4879] = ~(in[549] ^ in[521]); 
    assign layer_0[4880] = ~(in[262] ^ in[667]); 
    assign layer_0[4881] = 1'b1; 
    assign layer_0[4882] = ~(in[468] ^ in[355]); 
    assign layer_0[4883] = in[422] & ~in[266]; 
    assign layer_0[4884] = ~(in[239] & in[586]); 
    assign layer_0[4885] = ~in[552] | (in[552] & in[712]); 
    assign layer_0[4886] = ~in[340]; 
    assign layer_0[4887] = in[222] & ~in[275]; 
    assign layer_0[4888] = ~in[565] | (in[724] & in[565]); 
    assign layer_0[4889] = in[464] & ~in[154]; 
    assign layer_0[4890] = ~(in[39] ^ in[439]); 
    assign layer_0[4891] = in[388] ^ in[723]; 
    assign layer_0[4892] = ~(in[655] | in[42]); 
    assign layer_0[4893] = ~in[540]; 
    assign layer_0[4894] = ~(in[464] ^ in[312]); 
    assign layer_0[4895] = ~(in[97] ^ in[242]); 
    assign layer_0[4896] = in[424] ^ in[389]; 
    assign layer_0[4897] = ~(in[227] ^ in[598]); 
    assign layer_0[4898] = ~in[611]; 
    assign layer_0[4899] = in[6] | in[312]; 
    assign layer_0[4900] = in[294] & in[506]; 
    assign layer_0[4901] = in[439] & in[281]; 
    assign layer_0[4902] = in[47]; 
    assign layer_0[4903] = 1'b1; 
    assign layer_0[4904] = ~in[422] | (in[631] & in[422]); 
    assign layer_0[4905] = in[147] | in[532]; 
    assign layer_0[4906] = ~in[535] | (in[709] & in[535]); 
    assign layer_0[4907] = in[673] & ~in[69]; 
    assign layer_0[4908] = ~(in[185] | in[220]); 
    assign layer_0[4909] = in[276] ^ in[346]; 
    assign layer_0[4910] = ~(in[325] | in[331]); 
    assign layer_0[4911] = ~(in[205] & in[766]); 
    assign layer_0[4912] = ~(in[694] & in[409]); 
    assign layer_0[4913] = in[603] & ~in[552]; 
    assign layer_0[4914] = ~in[74] | (in[224] & in[74]); 
    assign layer_0[4915] = ~in[84] | (in[370] & in[84]); 
    assign layer_0[4916] = ~in[247]; 
    assign layer_0[4917] = ~(in[50] & in[379]); 
    assign layer_0[4918] = in[762] ^ in[650]; 
    assign layer_0[4919] = ~(in[395] & in[403]); 
    assign layer_0[4920] = ~(in[129] | in[452]); 
    assign layer_0[4921] = in[552]; 
    assign layer_0[4922] = ~(in[643] ^ in[325]); 
    assign layer_0[4923] = in[499] ^ in[464]; 
    assign layer_0[4924] = ~(in[372] ^ in[649]); 
    assign layer_0[4925] = ~(in[387] ^ in[380]); 
    assign layer_0[4926] = ~(in[30] & in[17]); 
    assign layer_0[4927] = 1'b1; 
    assign layer_0[4928] = in[595]; 
    assign layer_0[4929] = in[581] & ~in[651]; 
    assign layer_0[4930] = ~(in[653] | in[91]); 
    assign layer_0[4931] = in[435] & in[743]; 
    assign layer_0[4932] = ~in[50] | (in[246] & in[50]); 
    assign layer_0[4933] = ~(in[313] ^ in[504]); 
    assign layer_0[4934] = in[396] & ~in[138]; 
    assign layer_0[4935] = ~(in[371] ^ in[671]); 
    assign layer_0[4936] = ~(in[189] & in[479]); 
    assign layer_0[4937] = in[141] ^ in[648]; 
    assign layer_0[4938] = ~in[467]; 
    assign layer_0[4939] = ~(in[579] ^ in[412]); 
    assign layer_0[4940] = ~(in[324] & in[424]); 
    assign layer_0[4941] = in[311] ^ in[101]; 
    assign layer_0[4942] = in[538] | in[519]; 
    assign layer_0[4943] = ~in[360]; 
    assign layer_0[4944] = ~in[13] | (in[631] & in[13]); 
    assign layer_0[4945] = in[486] ^ in[265]; 
    assign layer_0[4946] = in[296] ^ in[724]; 
    assign layer_0[4947] = ~in[359] | (in[650] & in[359]); 
    assign layer_0[4948] = ~(in[659] ^ in[644]); 
    assign layer_0[4949] = in[739] & ~in[286]; 
    assign layer_0[4950] = ~in[194] | (in[289] & in[194]); 
    assign layer_0[4951] = ~in[671]; 
    assign layer_0[4952] = in[511] & ~in[492]; 
    assign layer_0[4953] = ~(in[684] | in[648]); 
    assign layer_0[4954] = ~in[703] | (in[703] & in[689]); 
    assign layer_0[4955] = in[213] ^ in[712]; 
    assign layer_0[4956] = ~(in[732] & in[551]); 
    assign layer_0[4957] = ~in[359] | (in[359] & in[699]); 
    assign layer_0[4958] = ~(in[106] ^ in[333]); 
    assign layer_0[4959] = in[186] | in[394]; 
    assign layer_0[4960] = ~in[220]; 
    assign layer_0[4961] = ~(in[504] | in[33]); 
    assign layer_0[4962] = in[147]; 
    assign layer_0[4963] = ~(in[502] ^ in[743]); 
    assign layer_0[4964] = ~(in[391] ^ in[489]); 
    assign layer_0[4965] = ~in[495]; 
    assign layer_0[4966] = in[403] & in[35]; 
    assign layer_0[4967] = ~(in[173] & in[205]); 
    assign layer_0[4968] = ~(in[701] ^ in[601]); 
    assign layer_0[4969] = in[469] & in[83]; 
    assign layer_0[4970] = in[325] | in[597]; 
    assign layer_0[4971] = ~in[582] | (in[597] & in[582]); 
    assign layer_0[4972] = ~in[328] | (in[647] & in[328]); 
    assign layer_0[4973] = ~in[24] | (in[24] & in[116]); 
    assign layer_0[4974] = ~(in[87] ^ in[417]); 
    assign layer_0[4975] = in[456] ^ in[36]; 
    assign layer_0[4976] = ~(in[84] & in[443]); 
    assign layer_0[4977] = in[309]; 
    assign layer_0[4978] = ~in[126]; 
    assign layer_0[4979] = in[741] ^ in[252]; 
    assign layer_0[4980] = in[349]; 
    assign layer_0[4981] = in[264] ^ in[266]; 
    assign layer_0[4982] = ~in[293]; 
    assign layer_0[4983] = in[343] ^ in[330]; 
    assign layer_0[4984] = ~(in[59] & in[428]); 
    assign layer_0[4985] = in[444] ^ in[127]; 
    assign layer_0[4986] = in[430]; 
    assign layer_0[4987] = in[263] ^ in[505]; 
    assign layer_0[4988] = in[4] & ~in[154]; 
    assign layer_0[4989] = in[187] & ~in[425]; 
    assign layer_0[4990] = in[649] & ~in[464]; 
    assign layer_0[4991] = in[280] & ~in[31]; 
    assign layer_0[4992] = ~(in[735] ^ in[623]); 
    assign layer_0[4993] = ~(in[713] ^ in[726]); 
    assign layer_0[4994] = ~(in[315] ^ in[518]); 
    assign layer_0[4995] = in[377]; 
    assign layer_0[4996] = in[575] & ~in[192]; 
    assign layer_0[4997] = ~in[340] | (in[191] & in[340]); 
    assign layer_0[4998] = ~in[762]; 
    assign layer_0[4999] = ~in[645] | (in[645] & in[12]); 
    assign layer_0[5000] = in[159] ^ in[8]; 
    assign layer_0[5001] = in[434] | in[79]; 
    assign layer_0[5002] = ~(in[696] ^ in[712]); 
    assign layer_0[5003] = in[7] & ~in[47]; 
    assign layer_0[5004] = in[663] & ~in[728]; 
    assign layer_0[5005] = ~in[530] | (in[435] & in[530]); 
    assign layer_0[5006] = in[81] ^ in[73]; 
    assign layer_0[5007] = ~in[321]; 
    assign layer_0[5008] = ~in[746] | (in[239] & in[746]); 
    assign layer_0[5009] = ~in[604]; 
    assign layer_0[5010] = in[109] & in[447]; 
    assign layer_0[5011] = ~(in[631] ^ in[3]); 
    assign layer_0[5012] = ~(in[627] ^ in[311]); 
    assign layer_0[5013] = ~in[204] | (in[204] & in[465]); 
    assign layer_0[5014] = ~(in[102] & in[571]); 
    assign layer_0[5015] = in[477] & in[254]; 
    assign layer_0[5016] = ~in[574]; 
    assign layer_0[5017] = ~(in[123] ^ in[601]); 
    assign layer_0[5018] = in[310] | in[337]; 
    assign layer_0[5019] = in[440] ^ in[422]; 
    assign layer_0[5020] = in[749]; 
    assign layer_0[5021] = ~in[174]; 
    assign layer_0[5022] = ~(in[602] ^ in[648]); 
    assign layer_0[5023] = in[226] & in[150]; 
    assign layer_0[5024] = in[458]; 
    assign layer_0[5025] = ~in[683]; 
    assign layer_0[5026] = in[684] | in[429]; 
    assign layer_0[5027] = in[47] ^ in[704]; 
    assign layer_0[5028] = in[491] ^ in[195]; 
    assign layer_0[5029] = in[344] & ~in[698]; 
    assign layer_0[5030] = in[11]; 
    assign layer_0[5031] = in[311]; 
    assign layer_0[5032] = ~in[419]; 
    assign layer_0[5033] = in[356] & ~in[744]; 
    assign layer_0[5034] = ~(in[445] & in[10]); 
    assign layer_0[5035] = ~in[494]; 
    assign layer_0[5036] = ~(in[282] ^ in[765]); 
    assign layer_0[5037] = ~in[654] | (in[654] & in[557]); 
    assign layer_0[5038] = ~in[331] | (in[360] & in[331]); 
    assign layer_0[5039] = in[387] ^ in[358]; 
    assign layer_0[5040] = in[229]; 
    assign layer_0[5041] = in[159]; 
    assign layer_0[5042] = ~(in[385] | in[468]); 
    assign layer_0[5043] = ~in[746]; 
    assign layer_0[5044] = in[261] ^ in[323]; 
    assign layer_0[5045] = ~in[462]; 
    assign layer_0[5046] = ~(in[553] ^ in[307]); 
    assign layer_0[5047] = ~(in[193] ^ in[452]); 
    assign layer_0[5048] = ~(in[474] ^ in[701]); 
    assign layer_0[5049] = ~(in[219] ^ in[17]); 
    assign layer_0[5050] = ~(in[300] & in[29]); 
    assign layer_0[5051] = in[468] & ~in[538]; 
    assign layer_0[5052] = ~in[731] | (in[731] & in[257]); 
    assign layer_0[5053] = ~(in[147] & in[265]); 
    assign layer_0[5054] = ~in[677] | (in[677] & in[673]); 
    assign layer_0[5055] = in[388] & ~in[196]; 
    assign layer_0[5056] = in[29]; 
    assign layer_0[5057] = ~in[52] | (in[61] & in[52]); 
    assign layer_0[5058] = in[265] & ~in[467]; 
    assign layer_0[5059] = ~in[594]; 
    assign layer_0[5060] = ~in[470] | (in[675] & in[470]); 
    assign layer_0[5061] = ~in[92]; 
    assign layer_0[5062] = ~in[518] | (in[244] & in[518]); 
    assign layer_0[5063] = in[3] ^ in[173]; 
    assign layer_0[5064] = ~(in[251] | in[632]); 
    assign layer_0[5065] = in[722] & ~in[260]; 
    assign layer_0[5066] = in[498] ^ in[542]; 
    assign layer_0[5067] = in[308] ^ in[551]; 
    assign layer_0[5068] = in[4]; 
    assign layer_0[5069] = ~in[25] | (in[25] & in[249]); 
    assign layer_0[5070] = ~(in[464] ^ in[437]); 
    assign layer_0[5071] = in[180] & ~in[530]; 
    assign layer_0[5072] = in[584] ^ in[666]; 
    assign layer_0[5073] = in[555]; 
    assign layer_0[5074] = in[403] | in[234]; 
    assign layer_0[5075] = in[338] ^ in[398]; 
    assign layer_0[5076] = in[636] ^ in[633]; 
    assign layer_0[5077] = ~(in[92] | in[28]); 
    assign layer_0[5078] = ~(in[290] ^ in[20]); 
    assign layer_0[5079] = ~in[536] | (in[536] & in[641]); 
    assign layer_0[5080] = ~in[647]; 
    assign layer_0[5081] = in[71] ^ in[52]; 
    assign layer_0[5082] = ~(in[466] ^ in[425]); 
    assign layer_0[5083] = in[633] ^ in[388]; 
    assign layer_0[5084] = in[634] | in[499]; 
    assign layer_0[5085] = in[182] & in[493]; 
    assign layer_0[5086] = ~in[457] | (in[457] & in[432]); 
    assign layer_0[5087] = in[601] ^ in[612]; 
    assign layer_0[5088] = in[334] ^ in[71]; 
    assign layer_0[5089] = in[633] & in[4]; 
    assign layer_0[5090] = in[553] ^ in[248]; 
    assign layer_0[5091] = in[352] | in[185]; 
    assign layer_0[5092] = ~in[583]; 
    assign layer_0[5093] = ~in[77] | (in[731] & in[77]); 
    assign layer_0[5094] = ~in[67]; 
    assign layer_0[5095] = ~in[747]; 
    assign layer_0[5096] = in[605]; 
    assign layer_0[5097] = ~(in[696] ^ in[697]); 
    assign layer_0[5098] = in[700] | in[450]; 
    assign layer_0[5099] = in[548]; 
    assign layer_0[5100] = ~(in[264] & in[440]); 
    assign layer_0[5101] = ~(in[467] ^ in[533]); 
    assign layer_0[5102] = ~in[27] | (in[282] & in[27]); 
    assign layer_0[5103] = in[145] & ~in[563]; 
    assign layer_0[5104] = in[19] & ~in[482]; 
    assign layer_0[5105] = in[599] & in[86]; 
    assign layer_0[5106] = ~in[8] | (in[8] & in[616]); 
    assign layer_0[5107] = ~(in[245] ^ in[448]); 
    assign layer_0[5108] = in[698]; 
    assign layer_0[5109] = in[453] & ~in[254]; 
    assign layer_0[5110] = in[717] ^ in[298]; 
    assign layer_0[5111] = ~(in[683] ^ in[190]); 
    assign layer_0[5112] = ~(in[500] ^ in[106]); 
    assign layer_0[5113] = in[294] & ~in[593]; 
    assign layer_0[5114] = ~(in[679] ^ in[680]); 
    assign layer_0[5115] = in[454] & in[346]; 
    assign layer_0[5116] = ~(in[148] ^ in[29]); 
    assign layer_0[5117] = in[459] & in[254]; 
    assign layer_0[5118] = ~in[490]; 
    assign layer_0[5119] = in[173] & ~in[476]; 
    assign layer_0[5120] = ~(in[302] & in[477]); 
    assign layer_0[5121] = ~in[81]; 
    assign layer_0[5122] = in[376] ^ in[380]; 
    assign layer_0[5123] = ~(in[420] ^ in[85]); 
    assign layer_0[5124] = in[329] ^ in[190]; 
    assign layer_0[5125] = in[230] ^ in[572]; 
    assign layer_0[5126] = in[507] ^ in[157]; 
    assign layer_0[5127] = in[456]; 
    assign layer_0[5128] = ~(in[724] | in[451]); 
    assign layer_0[5129] = ~(in[144] | in[284]); 
    assign layer_0[5130] = ~in[484] | (in[254] & in[484]); 
    assign layer_0[5131] = in[636] & ~in[599]; 
    assign layer_0[5132] = in[451] | in[379]; 
    assign layer_0[5133] = in[699] ^ in[412]; 
    assign layer_0[5134] = ~in[337]; 
    assign layer_0[5135] = ~in[291] | (in[291] & in[500]); 
    assign layer_0[5136] = ~in[501] | (in[34] & in[501]); 
    assign layer_0[5137] = in[538] ^ in[413]; 
    assign layer_0[5138] = ~(in[245] ^ in[572]); 
    assign layer_0[5139] = in[214] & in[4]; 
    assign layer_0[5140] = in[100] | in[17]; 
    assign layer_0[5141] = in[657]; 
    assign layer_0[5142] = in[341]; 
    assign layer_0[5143] = in[373] & in[606]; 
    assign layer_0[5144] = in[399] & ~in[682]; 
    assign layer_0[5145] = ~(in[553] | in[580]); 
    assign layer_0[5146] = in[728] & ~in[129]; 
    assign layer_0[5147] = in[61]; 
    assign layer_0[5148] = ~in[465] | (in[465] & in[544]); 
    assign layer_0[5149] = in[144] & ~in[736]; 
    assign layer_0[5150] = ~(in[553] ^ in[552]); 
    assign layer_0[5151] = in[362]; 
    assign layer_0[5152] = in[41]; 
    assign layer_0[5153] = ~(in[346] & in[376]); 
    assign layer_0[5154] = ~in[636]; 
    assign layer_0[5155] = ~(in[493] ^ in[430]); 
    assign layer_0[5156] = ~in[145]; 
    assign layer_0[5157] = ~in[613]; 
    assign layer_0[5158] = ~(in[331] & in[122]); 
    assign layer_0[5159] = in[689] & ~in[698]; 
    assign layer_0[5160] = in[425]; 
    assign layer_0[5161] = in[681] ^ in[374]; 
    assign layer_0[5162] = ~(in[292] | in[304]); 
    assign layer_0[5163] = ~(in[536] ^ in[565]); 
    assign layer_0[5164] = in[533] ^ in[210]; 
    assign layer_0[5165] = ~(in[462] & in[145]); 
    assign layer_0[5166] = ~in[567] | (in[567] & in[670]); 
    assign layer_0[5167] = in[659] & ~in[501]; 
    assign layer_0[5168] = in[325] & in[373]; 
    assign layer_0[5169] = 1'b0; 
    assign layer_0[5170] = in[251] ^ in[765]; 
    assign layer_0[5171] = ~(in[672] ^ in[416]); 
    assign layer_0[5172] = ~in[540]; 
    assign layer_0[5173] = in[141] | in[734]; 
    assign layer_0[5174] = in[660] ^ in[601]; 
    assign layer_0[5175] = in[709] | in[614]; 
    assign layer_0[5176] = in[393]; 
    assign layer_0[5177] = in[34] | in[130]; 
    assign layer_0[5178] = in[163] | in[219]; 
    assign layer_0[5179] = ~(in[450] ^ in[34]); 
    assign layer_0[5180] = in[664] ^ in[706]; 
    assign layer_0[5181] = ~in[252] | (in[370] & in[252]); 
    assign layer_0[5182] = in[537] | in[613]; 
    assign layer_0[5183] = in[654]; 
    assign layer_0[5184] = in[403] ^ in[586]; 
    assign layer_0[5185] = ~(in[11] ^ in[245]); 
    assign layer_0[5186] = ~in[68] | (in[68] & in[557]); 
    assign layer_0[5187] = ~in[180] | (in[339] & in[180]); 
    assign layer_0[5188] = ~in[535] | (in[535] & in[764]); 
    assign layer_0[5189] = ~in[129]; 
    assign layer_0[5190] = in[649] | in[733]; 
    assign layer_0[5191] = ~in[485]; 
    assign layer_0[5192] = ~(in[492] & in[196]); 
    assign layer_0[5193] = in[568]; 
    assign layer_0[5194] = ~in[455]; 
    assign layer_0[5195] = in[614] ^ in[720]; 
    assign layer_0[5196] = in[126] ^ in[373]; 
    assign layer_0[5197] = in[222] & ~in[506]; 
    assign layer_0[5198] = ~(in[615] ^ in[689]); 
    assign layer_0[5199] = ~in[81]; 
    assign layer_0[5200] = ~in[184]; 
    assign layer_0[5201] = in[691] & ~in[473]; 
    assign layer_0[5202] = in[236] & ~in[77]; 
    assign layer_0[5203] = in[264] & ~in[652]; 
    assign layer_0[5204] = ~(in[569] & in[237]); 
    assign layer_0[5205] = in[308] & ~in[531]; 
    assign layer_0[5206] = ~(in[689] ^ in[218]); 
    assign layer_0[5207] = ~in[472] | (in[519] & in[472]); 
    assign layer_0[5208] = ~(in[603] | in[62]); 
    assign layer_0[5209] = in[746]; 
    assign layer_0[5210] = in[61] ^ in[678]; 
    assign layer_0[5211] = in[234] & ~in[245]; 
    assign layer_0[5212] = in[394] & in[19]; 
    assign layer_0[5213] = in[598] & ~in[206]; 
    assign layer_0[5214] = ~in[67] | (in[67] & in[576]); 
    assign layer_0[5215] = in[549] ^ in[503]; 
    assign layer_0[5216] = ~in[742]; 
    assign layer_0[5217] = ~in[234] | (in[275] & in[234]); 
    assign layer_0[5218] = ~(in[174] ^ in[249]); 
    assign layer_0[5219] = in[575] & in[722]; 
    assign layer_0[5220] = in[712]; 
    assign layer_0[5221] = ~in[580] | (in[580] & in[501]); 
    assign layer_0[5222] = ~in[634]; 
    assign layer_0[5223] = in[378] & ~in[36]; 
    assign layer_0[5224] = ~(in[523] ^ in[716]); 
    assign layer_0[5225] = ~(in[435] | in[124]); 
    assign layer_0[5226] = ~(in[405] | in[209]); 
    assign layer_0[5227] = in[443] ^ in[746]; 
    assign layer_0[5228] = in[621] ^ in[579]; 
    assign layer_0[5229] = in[679]; 
    assign layer_0[5230] = in[98] & ~in[284]; 
    assign layer_0[5231] = in[177] & ~in[518]; 
    assign layer_0[5232] = ~in[146]; 
    assign layer_0[5233] = ~in[102]; 
    assign layer_0[5234] = ~(in[712] ^ in[424]); 
    assign layer_0[5235] = ~(in[245] & in[633]); 
    assign layer_0[5236] = in[253]; 
    assign layer_0[5237] = ~in[95] | (in[560] & in[95]); 
    assign layer_0[5238] = ~(in[681] ^ in[588]); 
    assign layer_0[5239] = ~in[735]; 
    assign layer_0[5240] = in[323] & in[759]; 
    assign layer_0[5241] = in[330]; 
    assign layer_0[5242] = in[650]; 
    assign layer_0[5243] = 1'b0; 
    assign layer_0[5244] = in[581] ^ in[20]; 
    assign layer_0[5245] = ~in[365]; 
    assign layer_0[5246] = ~in[381]; 
    assign layer_0[5247] = ~(in[78] ^ in[506]); 
    assign layer_0[5248] = ~(in[234] ^ in[102]); 
    assign layer_0[5249] = in[338] ^ in[680]; 
    assign layer_0[5250] = in[710] ^ in[712]; 
    assign layer_0[5251] = in[734] & ~in[410]; 
    assign layer_0[5252] = ~(in[656] ^ in[238]); 
    assign layer_0[5253] = in[413] & ~in[477]; 
    assign layer_0[5254] = ~(in[457] | in[609]); 
    assign layer_0[5255] = ~in[460] | (in[460] & in[630]); 
    assign layer_0[5256] = in[512] | in[357]; 
    assign layer_0[5257] = ~in[332] | (in[500] & in[332]); 
    assign layer_0[5258] = in[277] & in[506]; 
    assign layer_0[5259] = in[426] & ~in[229]; 
    assign layer_0[5260] = in[10] ^ in[426]; 
    assign layer_0[5261] = ~(in[108] ^ in[588]); 
    assign layer_0[5262] = in[23] | in[625]; 
    assign layer_0[5263] = in[201] ^ in[655]; 
    assign layer_0[5264] = in[756]; 
    assign layer_0[5265] = in[408] ^ in[730]; 
    assign layer_0[5266] = ~in[9]; 
    assign layer_0[5267] = ~(in[483] ^ in[619]); 
    assign layer_0[5268] = in[560] ^ in[363]; 
    assign layer_0[5269] = ~(in[729] & in[101]); 
    assign layer_0[5270] = in[404] | in[436]; 
    assign layer_0[5271] = ~in[520]; 
    assign layer_0[5272] = ~in[329]; 
    assign layer_0[5273] = in[585] ^ in[316]; 
    assign layer_0[5274] = in[631] | in[313]; 
    assign layer_0[5275] = in[652] & ~in[729]; 
    assign layer_0[5276] = ~(in[25] & in[440]); 
    assign layer_0[5277] = ~(in[683] ^ in[50]); 
    assign layer_0[5278] = ~(in[363] ^ in[520]); 
    assign layer_0[5279] = ~(in[694] ^ in[691]); 
    assign layer_0[5280] = ~(in[763] ^ in[680]); 
    assign layer_0[5281] = ~(in[416] ^ in[240]); 
    assign layer_0[5282] = ~in[255]; 
    assign layer_0[5283] = in[93] ^ in[246]; 
    assign layer_0[5284] = ~(in[282] & in[421]); 
    assign layer_0[5285] = ~in[98]; 
    assign layer_0[5286] = in[587] & in[82]; 
    assign layer_0[5287] = in[215] & ~in[302]; 
    assign layer_0[5288] = ~(in[392] & in[431]); 
    assign layer_0[5289] = in[53] & in[101]; 
    assign layer_0[5290] = in[572] ^ in[566]; 
    assign layer_0[5291] = in[300]; 
    assign layer_0[5292] = in[12]; 
    assign layer_0[5293] = ~in[238] | (in[605] & in[238]); 
    assign layer_0[5294] = ~in[428] | (in[579] & in[428]); 
    assign layer_0[5295] = in[195] & ~in[253]; 
    assign layer_0[5296] = in[283] ^ in[284]; 
    assign layer_0[5297] = ~in[664] | (in[758] & in[664]); 
    assign layer_0[5298] = in[246] & ~in[517]; 
    assign layer_0[5299] = ~(in[691] ^ in[728]); 
    assign layer_0[5300] = in[487] & in[520]; 
    assign layer_0[5301] = ~in[59] | (in[59] & in[284]); 
    assign layer_0[5302] = ~in[451]; 
    assign layer_0[5303] = in[317] ^ in[670]; 
    assign layer_0[5304] = in[559] | in[646]; 
    assign layer_0[5305] = ~(in[536] ^ in[339]); 
    assign layer_0[5306] = in[474] ^ in[339]; 
    assign layer_0[5307] = ~(in[676] ^ in[315]); 
    assign layer_0[5308] = ~(in[387] ^ in[494]); 
    assign layer_0[5309] = ~in[219]; 
    assign layer_0[5310] = in[1] ^ in[74]; 
    assign layer_0[5311] = in[12] & ~in[616]; 
    assign layer_0[5312] = in[262] & ~in[33]; 
    assign layer_0[5313] = in[73]; 
    assign layer_0[5314] = in[277] ^ in[250]; 
    assign layer_0[5315] = in[562] | in[1]; 
    assign layer_0[5316] = in[278] & ~in[651]; 
    assign layer_0[5317] = in[166] & ~in[461]; 
    assign layer_0[5318] = in[278] | in[294]; 
    assign layer_0[5319] = in[668] | in[65]; 
    assign layer_0[5320] = ~in[379]; 
    assign layer_0[5321] = ~in[645] | (in[645] & in[750]); 
    assign layer_0[5322] = ~(in[209] ^ in[567]); 
    assign layer_0[5323] = in[567] ^ in[343]; 
    assign layer_0[5324] = in[232]; 
    assign layer_0[5325] = ~(in[415] ^ in[399]); 
    assign layer_0[5326] = ~(in[601] ^ in[282]); 
    assign layer_0[5327] = in[514] & ~in[739]; 
    assign layer_0[5328] = in[332] & ~in[548]; 
    assign layer_0[5329] = in[202] ^ in[33]; 
    assign layer_0[5330] = ~(in[25] & in[122]); 
    assign layer_0[5331] = ~(in[622] & in[645]); 
    assign layer_0[5332] = in[525] ^ in[255]; 
    assign layer_0[5333] = ~(in[55] & in[27]); 
    assign layer_0[5334] = in[597] | in[16]; 
    assign layer_0[5335] = in[602]; 
    assign layer_0[5336] = ~(in[264] ^ in[260]); 
    assign layer_0[5337] = ~in[124] | (in[62] & in[124]); 
    assign layer_0[5338] = ~(in[342] & in[522]); 
    assign layer_0[5339] = in[372] & ~in[531]; 
    assign layer_0[5340] = ~in[98] | (in[98] & in[489]); 
    assign layer_0[5341] = ~(in[717] & in[469]); 
    assign layer_0[5342] = ~in[632] | (in[82] & in[632]); 
    assign layer_0[5343] = ~(in[266] & in[51]); 
    assign layer_0[5344] = in[461] ^ in[535]; 
    assign layer_0[5345] = ~in[392] | (in[204] & in[392]); 
    assign layer_0[5346] = in[348] & ~in[645]; 
    assign layer_0[5347] = in[679] ^ in[237]; 
    assign layer_0[5348] = ~in[396]; 
    assign layer_0[5349] = ~(in[647] ^ in[395]); 
    assign layer_0[5350] = ~(in[450] ^ in[716]); 
    assign layer_0[5351] = ~in[20]; 
    assign layer_0[5352] = ~(in[511] & in[52]); 
    assign layer_0[5353] = in[252] ^ in[586]; 
    assign layer_0[5354] = in[605] | in[14]; 
    assign layer_0[5355] = in[8] ^ in[753]; 
    assign layer_0[5356] = ~(in[75] ^ in[206]); 
    assign layer_0[5357] = ~in[65] | (in[65] & in[414]); 
    assign layer_0[5358] = ~(in[84] ^ in[570]); 
    assign layer_0[5359] = in[760] ^ in[759]; 
    assign layer_0[5360] = ~(in[293] ^ in[665]); 
    assign layer_0[5361] = ~(in[474] & in[472]); 
    assign layer_0[5362] = ~in[361] | (in[361] & in[598]); 
    assign layer_0[5363] = ~(in[698] ^ in[182]); 
    assign layer_0[5364] = in[404] ^ in[184]; 
    assign layer_0[5365] = ~in[716] | (in[716] & in[453]); 
    assign layer_0[5366] = ~in[250]; 
    assign layer_0[5367] = ~(in[460] ^ in[355]); 
    assign layer_0[5368] = in[448] ^ in[707]; 
    assign layer_0[5369] = in[464] & ~in[47]; 
    assign layer_0[5370] = ~(in[609] ^ in[737]); 
    assign layer_0[5371] = in[204] & ~in[396]; 
    assign layer_0[5372] = in[40] ^ in[728]; 
    assign layer_0[5373] = ~(in[93] & in[681]); 
    assign layer_0[5374] = ~in[607]; 
    assign layer_0[5375] = ~(in[666] ^ in[639]); 
    assign layer_0[5376] = ~(in[332] & in[298]); 
    assign layer_0[5377] = ~(in[177] ^ in[361]); 
    assign layer_0[5378] = ~(in[698] ^ in[501]); 
    assign layer_0[5379] = in[23] & in[112]; 
    assign layer_0[5380] = in[532] & in[422]; 
    assign layer_0[5381] = ~(in[232] ^ in[669]); 
    assign layer_0[5382] = ~in[455] | (in[482] & in[455]); 
    assign layer_0[5383] = ~in[262] | (in[262] & in[292]); 
    assign layer_0[5384] = in[217] & in[76]; 
    assign layer_0[5385] = in[590] & in[631]; 
    assign layer_0[5386] = in[396]; 
    assign layer_0[5387] = in[599] & ~in[604]; 
    assign layer_0[5388] = ~(in[568] ^ in[710]); 
    assign layer_0[5389] = ~(in[600] ^ in[620]); 
    assign layer_0[5390] = ~(in[300] ^ in[336]); 
    assign layer_0[5391] = ~(in[521] | in[762]); 
    assign layer_0[5392] = ~(in[673] | in[627]); 
    assign layer_0[5393] = ~(in[120] ^ in[402]); 
    assign layer_0[5394] = ~(in[254] ^ in[205]); 
    assign layer_0[5395] = in[730]; 
    assign layer_0[5396] = in[470]; 
    assign layer_0[5397] = in[348] & ~in[63]; 
    assign layer_0[5398] = in[582]; 
    assign layer_0[5399] = in[76] & ~in[704]; 
    assign layer_0[5400] = in[449]; 
    assign layer_0[5401] = ~(in[713] ^ in[66]); 
    assign layer_0[5402] = in[364] | in[310]; 
    assign layer_0[5403] = in[576] | in[642]; 
    assign layer_0[5404] = in[569] & in[695]; 
    assign layer_0[5405] = in[316] ^ in[670]; 
    assign layer_0[5406] = in[428] & in[537]; 
    assign layer_0[5407] = in[547] | in[673]; 
    assign layer_0[5408] = ~(in[341] ^ in[309]); 
    assign layer_0[5409] = in[521] ^ in[680]; 
    assign layer_0[5410] = ~(in[102] ^ in[275]); 
    assign layer_0[5411] = ~(in[669] ^ in[59]); 
    assign layer_0[5412] = in[473] | in[66]; 
    assign layer_0[5413] = ~(in[322] ^ in[265]); 
    assign layer_0[5414] = ~(in[322] & in[513]); 
    assign layer_0[5415] = in[2] & ~in[540]; 
    assign layer_0[5416] = in[530] ^ in[217]; 
    assign layer_0[5417] = in[581]; 
    assign layer_0[5418] = ~in[626]; 
    assign layer_0[5419] = in[666]; 
    assign layer_0[5420] = ~in[535] | (in[535] & in[541]); 
    assign layer_0[5421] = ~in[395] | (in[742] & in[395]); 
    assign layer_0[5422] = in[92] & ~in[49]; 
    assign layer_0[5423] = in[435] ^ in[707]; 
    assign layer_0[5424] = ~(in[111] & in[129]); 
    assign layer_0[5425] = in[716] ^ in[363]; 
    assign layer_0[5426] = ~in[644]; 
    assign layer_0[5427] = ~in[501] | (in[617] & in[501]); 
    assign layer_0[5428] = ~(in[424] ^ in[632]); 
    assign layer_0[5429] = ~(in[674] ^ in[70]); 
    assign layer_0[5430] = ~(in[267] ^ in[419]); 
    assign layer_0[5431] = in[162] ^ in[712]; 
    assign layer_0[5432] = in[593] | in[329]; 
    assign layer_0[5433] = in[344] ^ in[755]; 
    assign layer_0[5434] = in[373] & in[580]; 
    assign layer_0[5435] = in[28] ^ in[259]; 
    assign layer_0[5436] = in[446] ^ in[19]; 
    assign layer_0[5437] = ~in[665]; 
    assign layer_0[5438] = ~in[289]; 
    assign layer_0[5439] = ~(in[407] | in[664]); 
    assign layer_0[5440] = 1'b1; 
    assign layer_0[5441] = ~(in[259] | in[538]); 
    assign layer_0[5442] = in[341] & ~in[266]; 
    assign layer_0[5443] = ~(in[51] & in[628]); 
    assign layer_0[5444] = ~(in[583] ^ in[699]); 
    assign layer_0[5445] = in[388] & ~in[637]; 
    assign layer_0[5446] = in[501] & ~in[388]; 
    assign layer_0[5447] = ~(in[19] ^ in[661]); 
    assign layer_0[5448] = in[69] | in[630]; 
    assign layer_0[5449] = ~in[580] | (in[602] & in[580]); 
    assign layer_0[5450] = ~(in[142] ^ in[380]); 
    assign layer_0[5451] = ~(in[13] ^ in[146]); 
    assign layer_0[5452] = ~(in[589] | in[586]); 
    assign layer_0[5453] = in[399]; 
    assign layer_0[5454] = in[61]; 
    assign layer_0[5455] = ~in[341] | (in[341] & in[686]); 
    assign layer_0[5456] = in[674] | in[488]; 
    assign layer_0[5457] = ~(in[477] ^ in[660]); 
    assign layer_0[5458] = in[299] & ~in[468]; 
    assign layer_0[5459] = 1'b1; 
    assign layer_0[5460] = in[145] ^ in[646]; 
    assign layer_0[5461] = ~in[363] | (in[363] & in[1]); 
    assign layer_0[5462] = in[455] ^ in[454]; 
    assign layer_0[5463] = ~(in[21] & in[589]); 
    assign layer_0[5464] = ~(in[3] ^ in[584]); 
    assign layer_0[5465] = ~(in[636] ^ in[551]); 
    assign layer_0[5466] = ~in[465] | (in[465] & in[463]); 
    assign layer_0[5467] = ~(in[298] ^ in[748]); 
    assign layer_0[5468] = in[595]; 
    assign layer_0[5469] = ~(in[66] ^ in[476]); 
    assign layer_0[5470] = in[648] & in[654]; 
    assign layer_0[5471] = ~(in[174] ^ in[502]); 
    assign layer_0[5472] = ~(in[61] ^ in[679]); 
    assign layer_0[5473] = in[436] & ~in[741]; 
    assign layer_0[5474] = ~(in[219] | in[751]); 
    assign layer_0[5475] = in[10] & ~in[282]; 
    assign layer_0[5476] = in[619]; 
    assign layer_0[5477] = ~(in[193] ^ in[604]); 
    assign layer_0[5478] = ~(in[80] ^ in[336]); 
    assign layer_0[5479] = in[423] ^ in[212]; 
    assign layer_0[5480] = ~in[566] | (in[566] & in[586]); 
    assign layer_0[5481] = in[357] & ~in[493]; 
    assign layer_0[5482] = in[756] ^ in[513]; 
    assign layer_0[5483] = in[23] ^ in[86]; 
    assign layer_0[5484] = in[20]; 
    assign layer_0[5485] = in[629] & in[641]; 
    assign layer_0[5486] = ~(in[645] ^ in[698]); 
    assign layer_0[5487] = in[101] & ~in[79]; 
    assign layer_0[5488] = in[678] | in[184]; 
    assign layer_0[5489] = in[136] & ~in[66]; 
    assign layer_0[5490] = in[4] ^ in[401]; 
    assign layer_0[5491] = in[385] & ~in[298]; 
    assign layer_0[5492] = in[666]; 
    assign layer_0[5493] = ~in[291]; 
    assign layer_0[5494] = 1'b1; 
    assign layer_0[5495] = in[444] ^ in[252]; 
    assign layer_0[5496] = in[680] & ~in[309]; 
    assign layer_0[5497] = in[98] ^ in[8]; 
    assign layer_0[5498] = ~in[425]; 
    assign layer_0[5499] = ~(in[410] & in[644]); 
    assign layer_0[5500] = in[30] & in[745]; 
    assign layer_0[5501] = in[761] & ~in[268]; 
    assign layer_0[5502] = in[619] | in[529]; 
    assign layer_0[5503] = ~(in[245] ^ in[598]); 
    assign layer_0[5504] = in[454] & ~in[624]; 
    assign layer_0[5505] = in[59] & ~in[383]; 
    assign layer_0[5506] = ~(in[547] ^ in[445]); 
    assign layer_0[5507] = ~(in[340] | in[645]); 
    assign layer_0[5508] = ~in[261] | (in[15] & in[261]); 
    assign layer_0[5509] = in[289]; 
    assign layer_0[5510] = in[420] & ~in[47]; 
    assign layer_0[5511] = ~(in[464] | in[36]); 
    assign layer_0[5512] = in[326] ^ in[517]; 
    assign layer_0[5513] = in[652] ^ in[47]; 
    assign layer_0[5514] = ~in[43] | (in[739] & in[43]); 
    assign layer_0[5515] = in[484] | in[533]; 
    assign layer_0[5516] = in[627] ^ in[444]; 
    assign layer_0[5517] = ~in[662]; 
    assign layer_0[5518] = ~(in[710] | in[402]); 
    assign layer_0[5519] = ~(in[192] ^ in[386]); 
    assign layer_0[5520] = in[535] ^ in[533]; 
    assign layer_0[5521] = in[403]; 
    assign layer_0[5522] = 1'b0; 
    assign layer_0[5523] = in[637] ^ in[94]; 
    assign layer_0[5524] = ~(in[646] ^ in[628]); 
    assign layer_0[5525] = in[276] ^ in[708]; 
    assign layer_0[5526] = in[12] & in[27]; 
    assign layer_0[5527] = ~in[280] | (in[280] & in[364]); 
    assign layer_0[5528] = in[715] & ~in[567]; 
    assign layer_0[5529] = in[77]; 
    assign layer_0[5530] = in[177] ^ in[91]; 
    assign layer_0[5531] = ~(in[75] & in[587]); 
    assign layer_0[5532] = ~(in[361] ^ in[606]); 
    assign layer_0[5533] = in[614] & ~in[531]; 
    assign layer_0[5534] = ~(in[5] ^ in[338]); 
    assign layer_0[5535] = ~in[488] | (in[488] & in[357]); 
    assign layer_0[5536] = in[297]; 
    assign layer_0[5537] = ~(in[699] | in[732]); 
    assign layer_0[5538] = ~in[60] | (in[60] & in[701]); 
    assign layer_0[5539] = in[439] & ~in[1]; 
    assign layer_0[5540] = in[325]; 
    assign layer_0[5541] = in[698]; 
    assign layer_0[5542] = ~(in[677] ^ in[387]); 
    assign layer_0[5543] = in[459] ^ in[682]; 
    assign layer_0[5544] = ~(in[663] | in[477]); 
    assign layer_0[5545] = ~in[567] | (in[668] & in[567]); 
    assign layer_0[5546] = ~in[649]; 
    assign layer_0[5547] = in[568]; 
    assign layer_0[5548] = ~in[211] | (in[374] & in[211]); 
    assign layer_0[5549] = ~in[267]; 
    assign layer_0[5550] = ~in[661]; 
    assign layer_0[5551] = in[586] ^ in[603]; 
    assign layer_0[5552] = in[762] ^ in[519]; 
    assign layer_0[5553] = in[520]; 
    assign layer_0[5554] = ~in[602] | (in[599] & in[602]); 
    assign layer_0[5555] = ~in[397] | (in[397] & in[571]); 
    assign layer_0[5556] = in[53] | in[280]; 
    assign layer_0[5557] = in[326] ^ in[715]; 
    assign layer_0[5558] = ~(in[629] ^ in[728]); 
    assign layer_0[5559] = in[204] & ~in[506]; 
    assign layer_0[5560] = in[111] | in[751]; 
    assign layer_0[5561] = ~(in[307] | in[752]); 
    assign layer_0[5562] = in[57] & in[160]; 
    assign layer_0[5563] = ~in[349] | (in[756] & in[349]); 
    assign layer_0[5564] = in[664] | in[696]; 
    assign layer_0[5565] = ~(in[617] ^ in[554]); 
    assign layer_0[5566] = in[101] ^ in[192]; 
    assign layer_0[5567] = ~in[646]; 
    assign layer_0[5568] = ~(in[163] | in[492]); 
    assign layer_0[5569] = in[365]; 
    assign layer_0[5570] = in[485] | in[356]; 
    assign layer_0[5571] = in[489] & ~in[416]; 
    assign layer_0[5572] = in[396] & ~in[500]; 
    assign layer_0[5573] = in[633] ^ in[506]; 
    assign layer_0[5574] = in[548] | in[660]; 
    assign layer_0[5575] = in[270]; 
    assign layer_0[5576] = in[587] & in[630]; 
    assign layer_0[5577] = ~(in[379] ^ in[499]); 
    assign layer_0[5578] = ~(in[501] ^ in[97]); 
    assign layer_0[5579] = in[51] & ~in[537]; 
    assign layer_0[5580] = ~in[743] | (in[743] & in[650]); 
    assign layer_0[5581] = in[597] & ~in[457]; 
    assign layer_0[5582] = in[739] | in[311]; 
    assign layer_0[5583] = in[394] & in[634]; 
    assign layer_0[5584] = ~(in[756] ^ in[615]); 
    assign layer_0[5585] = in[8]; 
    assign layer_0[5586] = ~in[416]; 
    assign layer_0[5587] = in[489] & in[180]; 
    assign layer_0[5588] = in[587] ^ in[583]; 
    assign layer_0[5589] = ~in[728]; 
    assign layer_0[5590] = ~(in[681] | in[11]); 
    assign layer_0[5591] = ~(in[650] ^ in[78]); 
    assign layer_0[5592] = ~(in[193] ^ in[292]); 
    assign layer_0[5593] = ~(in[69] ^ in[334]); 
    assign layer_0[5594] = in[362] & ~in[627]; 
    assign layer_0[5595] = in[507] ^ in[456]; 
    assign layer_0[5596] = in[699] & in[392]; 
    assign layer_0[5597] = in[295] & ~in[45]; 
    assign layer_0[5598] = ~in[376] | (in[360] & in[376]); 
    assign layer_0[5599] = in[596] ^ in[149]; 
    assign layer_0[5600] = ~(in[731] ^ in[326]); 
    assign layer_0[5601] = ~(in[348] & in[365]); 
    assign layer_0[5602] = in[296] | in[612]; 
    assign layer_0[5603] = ~in[656] | (in[656] & in[293]); 
    assign layer_0[5604] = in[374] & ~in[491]; 
    assign layer_0[5605] = ~(in[66] ^ in[62]); 
    assign layer_0[5606] = ~(in[599] & in[131]); 
    assign layer_0[5607] = in[291] | in[145]; 
    assign layer_0[5608] = ~in[458] | (in[458] & in[760]); 
    assign layer_0[5609] = ~in[312] | (in[312] & in[536]); 
    assign layer_0[5610] = in[283] ^ in[507]; 
    assign layer_0[5611] = in[731] ^ in[437]; 
    assign layer_0[5612] = in[315]; 
    assign layer_0[5613] = ~in[348] | (in[18] & in[348]); 
    assign layer_0[5614] = ~(in[69] ^ in[638]); 
    assign layer_0[5615] = in[658] | in[27]; 
    assign layer_0[5616] = ~(in[606] ^ in[659]); 
    assign layer_0[5617] = in[348]; 
    assign layer_0[5618] = in[50] & ~in[436]; 
    assign layer_0[5619] = in[708] & ~in[585]; 
    assign layer_0[5620] = in[367]; 
    assign layer_0[5621] = ~(in[292] ^ in[249]); 
    assign layer_0[5622] = in[277] ^ in[364]; 
    assign layer_0[5623] = ~in[641] | (in[641] & in[463]); 
    assign layer_0[5624] = ~in[714] | (in[714] & in[633]); 
    assign layer_0[5625] = in[37]; 
    assign layer_0[5626] = ~in[166]; 
    assign layer_0[5627] = in[604] ^ in[78]; 
    assign layer_0[5628] = ~in[426] | (in[426] & in[624]); 
    assign layer_0[5629] = ~(in[211] ^ in[710]); 
    assign layer_0[5630] = in[292]; 
    assign layer_0[5631] = ~(in[659] | in[227]); 
    assign layer_0[5632] = ~in[239]; 
    assign layer_0[5633] = ~in[411]; 
    assign layer_0[5634] = in[101]; 
    assign layer_0[5635] = ~(in[126] ^ in[597]); 
    assign layer_0[5636] = in[314] & ~in[693]; 
    assign layer_0[5637] = ~in[509] | (in[760] & in[509]); 
    assign layer_0[5638] = ~in[307]; 
    assign layer_0[5639] = in[503] & ~in[699]; 
    assign layer_0[5640] = in[679] ^ in[110]; 
    assign layer_0[5641] = in[102] ^ in[417]; 
    assign layer_0[5642] = in[154] & ~in[356]; 
    assign layer_0[5643] = ~(in[100] ^ in[673]); 
    assign layer_0[5644] = in[143] & ~in[704]; 
    assign layer_0[5645] = in[707] | in[220]; 
    assign layer_0[5646] = in[196]; 
    assign layer_0[5647] = in[37] & in[188]; 
    assign layer_0[5648] = ~(in[153] & in[391]); 
    assign layer_0[5649] = in[316] ^ in[504]; 
    assign layer_0[5650] = ~(in[437] ^ in[739]); 
    assign layer_0[5651] = in[8] | in[276]; 
    assign layer_0[5652] = in[263]; 
    assign layer_0[5653] = in[727] ^ in[635]; 
    assign layer_0[5654] = in[356] & ~in[520]; 
    assign layer_0[5655] = in[564] & ~in[701]; 
    assign layer_0[5656] = in[499]; 
    assign layer_0[5657] = in[579] ^ in[666]; 
    assign layer_0[5658] = in[84]; 
    assign layer_0[5659] = ~in[476]; 
    assign layer_0[5660] = in[570] ^ in[634]; 
    assign layer_0[5661] = in[272] ^ in[20]; 
    assign layer_0[5662] = ~(in[632] | in[232]); 
    assign layer_0[5663] = in[211] ^ in[340]; 
    assign layer_0[5664] = in[478] | in[288]; 
    assign layer_0[5665] = ~in[330]; 
    assign layer_0[5666] = ~in[578] | (in[578] & in[518]); 
    assign layer_0[5667] = in[9] & ~in[316]; 
    assign layer_0[5668] = in[358] ^ in[742]; 
    assign layer_0[5669] = ~(in[631] | in[658]); 
    assign layer_0[5670] = ~in[17]; 
    assign layer_0[5671] = ~(in[666] ^ in[458]); 
    assign layer_0[5672] = ~in[118] | (in[304] & in[118]); 
    assign layer_0[5673] = in[217] & in[727]; 
    assign layer_0[5674] = ~(in[486] ^ in[627]); 
    assign layer_0[5675] = ~in[237] | (in[237] & in[502]); 
    assign layer_0[5676] = ~(in[638] ^ in[94]); 
    assign layer_0[5677] = ~(in[339] | in[586]); 
    assign layer_0[5678] = 1'b0; 
    assign layer_0[5679] = in[347] ^ in[426]; 
    assign layer_0[5680] = ~in[252] | (in[725] & in[252]); 
    assign layer_0[5681] = in[79] ^ in[727]; 
    assign layer_0[5682] = in[294] | in[657]; 
    assign layer_0[5683] = ~(in[534] ^ in[569]); 
    assign layer_0[5684] = in[506] & ~in[34]; 
    assign layer_0[5685] = in[762]; 
    assign layer_0[5686] = in[647] & ~in[754]; 
    assign layer_0[5687] = in[598] ^ in[574]; 
    assign layer_0[5688] = in[235] | in[322]; 
    assign layer_0[5689] = ~(in[745] | in[365]); 
    assign layer_0[5690] = ~(in[88] ^ in[705]); 
    assign layer_0[5691] = in[611] ^ in[646]; 
    assign layer_0[5692] = ~in[347]; 
    assign layer_0[5693] = ~in[80]; 
    assign layer_0[5694] = in[690] ^ in[299]; 
    assign layer_0[5695] = in[427] & in[179]; 
    assign layer_0[5696] = in[348] & in[603]; 
    assign layer_0[5697] = ~in[660] | (in[660] & in[440]); 
    assign layer_0[5698] = ~(in[639] ^ in[613]); 
    assign layer_0[5699] = in[711]; 
    assign layer_0[5700] = in[744]; 
    assign layer_0[5701] = in[644] ^ in[621]; 
    assign layer_0[5702] = ~(in[567] ^ in[283]); 
    assign layer_0[5703] = in[629] | in[612]; 
    assign layer_0[5704] = in[361] ^ in[553]; 
    assign layer_0[5705] = ~in[53]; 
    assign layer_0[5706] = ~(in[344] ^ in[66]); 
    assign layer_0[5707] = in[693] & in[288]; 
    assign layer_0[5708] = in[659] ^ in[38]; 
    assign layer_0[5709] = in[720]; 
    assign layer_0[5710] = ~(in[287] | in[65]); 
    assign layer_0[5711] = ~(in[90] ^ in[604]); 
    assign layer_0[5712] = ~(in[618] & in[614]); 
    assign layer_0[5713] = ~in[51] | (in[51] & in[550]); 
    assign layer_0[5714] = ~(in[619] ^ in[370]); 
    assign layer_0[5715] = ~in[111] | (in[480] & in[111]); 
    assign layer_0[5716] = in[492] & ~in[701]; 
    assign layer_0[5717] = 1'b1; 
    assign layer_0[5718] = ~in[453]; 
    assign layer_0[5719] = ~(in[72] ^ in[417]); 
    assign layer_0[5720] = in[357] & ~in[689]; 
    assign layer_0[5721] = in[518] ^ in[344]; 
    assign layer_0[5722] = ~in[664]; 
    assign layer_0[5723] = in[659]; 
    assign layer_0[5724] = in[678] ^ in[519]; 
    assign layer_0[5725] = in[169] ^ in[519]; 
    assign layer_0[5726] = in[638] & in[349]; 
    assign layer_0[5727] = ~in[587]; 
    assign layer_0[5728] = in[428] | in[19]; 
    assign layer_0[5729] = in[592] | in[210]; 
    assign layer_0[5730] = ~(in[696] & in[670]); 
    assign layer_0[5731] = ~(in[514] ^ in[667]); 
    assign layer_0[5732] = ~in[606]; 
    assign layer_0[5733] = ~in[99] | (in[95] & in[99]); 
    assign layer_0[5734] = ~in[762] | (in[669] & in[762]); 
    assign layer_0[5735] = in[391] & in[476]; 
    assign layer_0[5736] = ~in[115] | (in[115] & in[707]); 
    assign layer_0[5737] = in[310] ^ in[614]; 
    assign layer_0[5738] = ~in[699] | (in[699] & in[601]); 
    assign layer_0[5739] = in[312]; 
    assign layer_0[5740] = in[685] ^ in[743]; 
    assign layer_0[5741] = ~(in[747] | in[264]); 
    assign layer_0[5742] = in[462] ^ in[78]; 
    assign layer_0[5743] = in[579] ^ in[355]; 
    assign layer_0[5744] = ~in[455] | (in[455] & in[93]); 
    assign layer_0[5745] = in[417] ^ in[278]; 
    assign layer_0[5746] = in[611] & in[393]; 
    assign layer_0[5747] = in[695] & ~in[380]; 
    assign layer_0[5748] = ~(in[34] | in[145]); 
    assign layer_0[5749] = ~in[184]; 
    assign layer_0[5750] = in[741]; 
    assign layer_0[5751] = in[89] & ~in[337]; 
    assign layer_0[5752] = ~in[25]; 
    assign layer_0[5753] = ~in[428]; 
    assign layer_0[5754] = ~in[357]; 
    assign layer_0[5755] = in[607] ^ in[200]; 
    assign layer_0[5756] = in[27]; 
    assign layer_0[5757] = ~(in[492] | in[700]); 
    assign layer_0[5758] = in[326] & ~in[595]; 
    assign layer_0[5759] = ~(in[462] | in[116]); 
    assign layer_0[5760] = in[500] ^ in[277]; 
    assign layer_0[5761] = in[332] & in[244]; 
    assign layer_0[5762] = in[5] & ~in[563]; 
    assign layer_0[5763] = in[311] & ~in[29]; 
    assign layer_0[5764] = ~(in[586] ^ in[628]); 
    assign layer_0[5765] = ~(in[659] ^ in[360]); 
    assign layer_0[5766] = in[576]; 
    assign layer_0[5767] = ~(in[584] ^ in[645]); 
    assign layer_0[5768] = ~(in[674] | in[767]); 
    assign layer_0[5769] = ~in[443] | (in[395] & in[443]); 
    assign layer_0[5770] = in[554] & ~in[636]; 
    assign layer_0[5771] = in[448]; 
    assign layer_0[5772] = in[656] ^ in[518]; 
    assign layer_0[5773] = ~(in[507] ^ in[205]); 
    assign layer_0[5774] = ~in[172]; 
    assign layer_0[5775] = in[113] ^ in[602]; 
    assign layer_0[5776] = ~in[574]; 
    assign layer_0[5777] = in[319] | in[329]; 
    assign layer_0[5778] = in[451] & ~in[664]; 
    assign layer_0[5779] = ~in[324]; 
    assign layer_0[5780] = ~(in[554] | in[598]); 
    assign layer_0[5781] = in[255] | in[400]; 
    assign layer_0[5782] = ~(in[357] ^ in[617]); 
    assign layer_0[5783] = ~in[424] | (in[424] & in[701]); 
    assign layer_0[5784] = ~in[753] | (in[21] & in[753]); 
    assign layer_0[5785] = in[380] & in[598]; 
    assign layer_0[5786] = ~(in[533] ^ in[281]); 
    assign layer_0[5787] = ~(in[192] ^ in[393]); 
    assign layer_0[5788] = in[298] & ~in[365]; 
    assign layer_0[5789] = ~(in[532] ^ in[328]); 
    assign layer_0[5790] = ~in[538] | (in[435] & in[538]); 
    assign layer_0[5791] = in[632] ^ in[630]; 
    assign layer_0[5792] = ~(in[34] ^ in[453]); 
    assign layer_0[5793] = in[469]; 
    assign layer_0[5794] = in[641] ^ in[697]; 
    assign layer_0[5795] = ~(in[525] | in[337]); 
    assign layer_0[5796] = ~in[88] | (in[319] & in[88]); 
    assign layer_0[5797] = ~in[451] | (in[451] & in[759]); 
    assign layer_0[5798] = in[156] & ~in[300]; 
    assign layer_0[5799] = ~(in[309] ^ in[123]); 
    assign layer_0[5800] = in[725] ^ in[147]; 
    assign layer_0[5801] = ~(in[679] ^ in[499]); 
    assign layer_0[5802] = in[633] ^ in[622]; 
    assign layer_0[5803] = ~in[10]; 
    assign layer_0[5804] = in[222] & ~in[303]; 
    assign layer_0[5805] = ~(in[451] | in[460]); 
    assign layer_0[5806] = ~(in[535] ^ in[556]); 
    assign layer_0[5807] = in[551] ^ in[316]; 
    assign layer_0[5808] = in[564] & in[387]; 
    assign layer_0[5809] = in[470] ^ in[48]; 
    assign layer_0[5810] = in[631] ^ in[569]; 
    assign layer_0[5811] = in[519]; 
    assign layer_0[5812] = in[173]; 
    assign layer_0[5813] = in[127]; 
    assign layer_0[5814] = in[660] ^ in[763]; 
    assign layer_0[5815] = ~in[673] | (in[311] & in[673]); 
    assign layer_0[5816] = ~(in[743] ^ in[178]); 
    assign layer_0[5817] = ~in[475]; 
    assign layer_0[5818] = ~in[421]; 
    assign layer_0[5819] = ~(in[269] | in[510]); 
    assign layer_0[5820] = ~in[452]; 
    assign layer_0[5821] = in[641]; 
    assign layer_0[5822] = in[224] ^ in[757]; 
    assign layer_0[5823] = in[284]; 
    assign layer_0[5824] = ~(in[580] ^ in[142]); 
    assign layer_0[5825] = ~(in[573] | in[239]); 
    assign layer_0[5826] = in[133]; 
    assign layer_0[5827] = in[286] | in[679]; 
    assign layer_0[5828] = ~(in[614] & in[312]); 
    assign layer_0[5829] = ~(in[605] | in[267]); 
    assign layer_0[5830] = in[711] & in[265]; 
    assign layer_0[5831] = in[60] ^ in[405]; 
    assign layer_0[5832] = in[304] | in[260]; 
    assign layer_0[5833] = in[689] & ~in[466]; 
    assign layer_0[5834] = ~in[68]; 
    assign layer_0[5835] = ~(in[587] | in[573]); 
    assign layer_0[5836] = ~(in[65] & in[64]); 
    assign layer_0[5837] = ~(in[571] ^ in[266]); 
    assign layer_0[5838] = ~in[401]; 
    assign layer_0[5839] = ~(in[324] ^ in[566]); 
    assign layer_0[5840] = ~in[323]; 
    assign layer_0[5841] = in[331] & ~in[413]; 
    assign layer_0[5842] = ~(in[573] | in[386]); 
    assign layer_0[5843] = in[476] | in[157]; 
    assign layer_0[5844] = ~(in[333] ^ in[388]); 
    assign layer_0[5845] = ~(in[596] | in[443]); 
    assign layer_0[5846] = ~in[143]; 
    assign layer_0[5847] = in[759] ^ in[677]; 
    assign layer_0[5848] = ~(in[646] ^ in[60]); 
    assign layer_0[5849] = ~(in[588] ^ in[253]); 
    assign layer_0[5850] = ~(in[186] & in[660]); 
    assign layer_0[5851] = ~in[234] | (in[413] & in[234]); 
    assign layer_0[5852] = ~(in[13] ^ in[446]); 
    assign layer_0[5853] = in[691] & ~in[282]; 
    assign layer_0[5854] = in[277] & ~in[264]; 
    assign layer_0[5855] = in[260] | in[552]; 
    assign layer_0[5856] = ~(in[667] | in[370]); 
    assign layer_0[5857] = ~(in[56] & in[731]); 
    assign layer_0[5858] = 1'b1; 
    assign layer_0[5859] = ~in[118] | (in[628] & in[118]); 
    assign layer_0[5860] = ~(in[62] ^ in[457]); 
    assign layer_0[5861] = in[104] & in[13]; 
    assign layer_0[5862] = ~(in[439] ^ in[391]); 
    assign layer_0[5863] = in[88] & ~in[137]; 
    assign layer_0[5864] = ~in[649]; 
    assign layer_0[5865] = ~(in[687] ^ in[432]); 
    assign layer_0[5866] = in[140]; 
    assign layer_0[5867] = in[505]; 
    assign layer_0[5868] = in[744] | in[159]; 
    assign layer_0[5869] = ~in[478]; 
    assign layer_0[5870] = in[730] ^ in[332]; 
    assign layer_0[5871] = in[329] | in[511]; 
    assign layer_0[5872] = in[614] ^ in[602]; 
    assign layer_0[5873] = ~in[520] | (in[84] & in[520]); 
    assign layer_0[5874] = ~(in[301] & in[714]); 
    assign layer_0[5875] = in[592] & ~in[333]; 
    assign layer_0[5876] = ~in[536] | (in[300] & in[536]); 
    assign layer_0[5877] = ~in[679]; 
    assign layer_0[5878] = ~(in[70] & in[125]); 
    assign layer_0[5879] = ~(in[498] & in[617]); 
    assign layer_0[5880] = in[676] ^ in[75]; 
    assign layer_0[5881] = ~(in[172] ^ in[73]); 
    assign layer_0[5882] = in[639]; 
    assign layer_0[5883] = ~in[147] | (in[668] & in[147]); 
    assign layer_0[5884] = in[251]; 
    assign layer_0[5885] = ~(in[579] & in[274]); 
    assign layer_0[5886] = in[502] | in[718]; 
    assign layer_0[5887] = ~in[455] | (in[455] & in[225]); 
    assign layer_0[5888] = in[633] | in[491]; 
    assign layer_0[5889] = in[584] & in[145]; 
    assign layer_0[5890] = in[726] ^ in[137]; 
    assign layer_0[5891] = ~in[5]; 
    assign layer_0[5892] = in[718] ^ in[493]; 
    assign layer_0[5893] = ~(in[212] | in[437]); 
    assign layer_0[5894] = in[68] ^ in[550]; 
    assign layer_0[5895] = in[477]; 
    assign layer_0[5896] = in[103] & in[344]; 
    assign layer_0[5897] = in[549] ^ in[10]; 
    assign layer_0[5898] = in[396] & ~in[110]; 
    assign layer_0[5899] = ~(in[61] ^ in[3]); 
    assign layer_0[5900] = in[230] & ~in[2]; 
    assign layer_0[5901] = in[729]; 
    assign layer_0[5902] = in[740] ^ in[604]; 
    assign layer_0[5903] = ~(in[417] ^ in[299]); 
    assign layer_0[5904] = in[707] ^ in[396]; 
    assign layer_0[5905] = ~in[385]; 
    assign layer_0[5906] = ~(in[516] | in[740]); 
    assign layer_0[5907] = in[619] ^ in[648]; 
    assign layer_0[5908] = ~in[485] | (in[590] & in[485]); 
    assign layer_0[5909] = in[107] ^ in[299]; 
    assign layer_0[5910] = in[396] ^ in[548]; 
    assign layer_0[5911] = in[94] ^ in[405]; 
    assign layer_0[5912] = ~in[429]; 
    assign layer_0[5913] = in[467] ^ in[93]; 
    assign layer_0[5914] = ~(in[616] ^ in[701]); 
    assign layer_0[5915] = ~in[324] | (in[324] & in[518]); 
    assign layer_0[5916] = in[253] ^ in[632]; 
    assign layer_0[5917] = in[628] & ~in[467]; 
    assign layer_0[5918] = in[292] & ~in[459]; 
    assign layer_0[5919] = in[486] & in[765]; 
    assign layer_0[5920] = ~(in[737] | in[330]); 
    assign layer_0[5921] = in[83] & in[314]; 
    assign layer_0[5922] = ~(in[725] & in[757]); 
    assign layer_0[5923] = ~(in[307] ^ in[453]); 
    assign layer_0[5924] = in[597] ^ in[434]; 
    assign layer_0[5925] = ~in[350] | (in[297] & in[350]); 
    assign layer_0[5926] = ~(in[5] & in[474]); 
    assign layer_0[5927] = in[239] ^ in[207]; 
    assign layer_0[5928] = ~in[370]; 
    assign layer_0[5929] = ~(in[739] & in[435]); 
    assign layer_0[5930] = in[279] ^ in[396]; 
    assign layer_0[5931] = ~(in[466] ^ in[468]); 
    assign layer_0[5932] = in[762] ^ in[232]; 
    assign layer_0[5933] = in[208] ^ in[385]; 
    assign layer_0[5934] = ~(in[260] ^ in[141]); 
    assign layer_0[5935] = ~(in[242] & in[253]); 
    assign layer_0[5936] = ~in[61] | (in[752] & in[61]); 
    assign layer_0[5937] = ~in[349] | (in[349] & in[191]); 
    assign layer_0[5938] = ~in[377]; 
    assign layer_0[5939] = in[315] ^ in[476]; 
    assign layer_0[5940] = in[648] & in[418]; 
    assign layer_0[5941] = in[261] ^ in[563]; 
    assign layer_0[5942] = in[654] & ~in[221]; 
    assign layer_0[5943] = ~in[632]; 
    assign layer_0[5944] = in[370]; 
    assign layer_0[5945] = ~in[160] | (in[160] & in[400]); 
    assign layer_0[5946] = in[319] | in[727]; 
    assign layer_0[5947] = ~in[682]; 
    assign layer_0[5948] = ~(in[205] ^ in[661]); 
    assign layer_0[5949] = in[218] & in[226]; 
    assign layer_0[5950] = in[552] & in[668]; 
    assign layer_0[5951] = in[650] | in[619]; 
    assign layer_0[5952] = ~in[537] | (in[537] & in[274]); 
    assign layer_0[5953] = in[449] ^ in[689]; 
    assign layer_0[5954] = ~(in[715] ^ in[670]); 
    assign layer_0[5955] = in[488] & ~in[743]; 
    assign layer_0[5956] = in[718]; 
    assign layer_0[5957] = ~in[78] | (in[78] & in[494]); 
    assign layer_0[5958] = ~in[50] | (in[50] & in[248]); 
    assign layer_0[5959] = in[555] ^ in[514]; 
    assign layer_0[5960] = in[371] | in[480]; 
    assign layer_0[5961] = in[333] | in[242]; 
    assign layer_0[5962] = in[326] & ~in[605]; 
    assign layer_0[5963] = in[709] & in[715]; 
    assign layer_0[5964] = ~(in[253] & in[277]); 
    assign layer_0[5965] = ~in[20] | (in[20] & in[642]); 
    assign layer_0[5966] = in[519] ^ in[518]; 
    assign layer_0[5967] = in[262] & ~in[178]; 
    assign layer_0[5968] = in[83] | in[704]; 
    assign layer_0[5969] = ~(in[388] & in[458]); 
    assign layer_0[5970] = ~in[600]; 
    assign layer_0[5971] = ~(in[211] ^ in[241]); 
    assign layer_0[5972] = in[674] ^ in[478]; 
    assign layer_0[5973] = in[604] & ~in[257]; 
    assign layer_0[5974] = in[187] & ~in[283]; 
    assign layer_0[5975] = in[3]; 
    assign layer_0[5976] = ~in[372]; 
    assign layer_0[5977] = in[333] & in[292]; 
    assign layer_0[5978] = in[538]; 
    assign layer_0[5979] = ~(in[279] & in[501]); 
    assign layer_0[5980] = ~in[322]; 
    assign layer_0[5981] = ~(in[509] | in[597]); 
    assign layer_0[5982] = in[451] & ~in[20]; 
    assign layer_0[5983] = in[659] ^ in[694]; 
    assign layer_0[5984] = in[636] | in[656]; 
    assign layer_0[5985] = ~in[164]; 
    assign layer_0[5986] = ~in[28]; 
    assign layer_0[5987] = in[533] & ~in[236]; 
    assign layer_0[5988] = in[454] & ~in[300]; 
    assign layer_0[5989] = ~in[384] | (in[217] & in[384]); 
    assign layer_0[5990] = ~(in[211] & in[105]); 
    assign layer_0[5991] = in[56] & ~in[209]; 
    assign layer_0[5992] = in[568] & ~in[35]; 
    assign layer_0[5993] = ~in[394] | (in[394] & in[631]); 
    assign layer_0[5994] = in[141] ^ in[380]; 
    assign layer_0[5995] = in[106] & ~in[460]; 
    assign layer_0[5996] = ~in[162] | (in[581] & in[162]); 
    assign layer_0[5997] = in[181] & in[122]; 
    assign layer_0[5998] = ~in[12]; 
    assign layer_0[5999] = in[205] ^ in[173]; 
    assign layer_0[6000] = in[333] | in[469]; 
    assign layer_0[6001] = ~in[208]; 
    assign layer_0[6002] = ~(in[648] ^ in[650]); 
    assign layer_0[6003] = in[471] & ~in[246]; 
    assign layer_0[6004] = in[11]; 
    assign layer_0[6005] = in[724] & in[494]; 
    assign layer_0[6006] = in[378] ^ in[424]; 
    assign layer_0[6007] = in[428] & ~in[673]; 
    assign layer_0[6008] = in[266] ^ in[410]; 
    assign layer_0[6009] = in[429] & ~in[249]; 
    assign layer_0[6010] = in[455] & ~in[365]; 
    assign layer_0[6011] = ~(in[723] ^ in[248]); 
    assign layer_0[6012] = in[476] ^ in[92]; 
    assign layer_0[6013] = ~in[710] | (in[714] & in[710]); 
    assign layer_0[6014] = in[187] | in[724]; 
    assign layer_0[6015] = in[307]; 
    assign layer_0[6016] = in[595] ^ in[759]; 
    assign layer_0[6017] = ~(in[169] ^ in[212]); 
    assign layer_0[6018] = ~in[438] | (in[438] & in[418]); 
    assign layer_0[6019] = in[694] ^ in[729]; 
    assign layer_0[6020] = ~(in[346] | in[336]); 
    assign layer_0[6021] = in[636] ^ in[4]; 
    assign layer_0[6022] = ~in[63] | (in[63] & in[133]); 
    assign layer_0[6023] = ~in[427]; 
    assign layer_0[6024] = in[649] ^ in[568]; 
    assign layer_0[6025] = in[264] & in[485]; 
    assign layer_0[6026] = in[471]; 
    assign layer_0[6027] = in[662] ^ in[476]; 
    assign layer_0[6028] = in[677] & ~in[602]; 
    assign layer_0[6029] = ~(in[244] ^ in[444]); 
    assign layer_0[6030] = ~in[78]; 
    assign layer_0[6031] = in[740] ^ in[83]; 
    assign layer_0[6032] = ~in[647]; 
    assign layer_0[6033] = ~(in[726] ^ in[725]); 
    assign layer_0[6034] = in[479] ^ in[311]; 
    assign layer_0[6035] = ~(in[579] & in[650]); 
    assign layer_0[6036] = in[432] ^ in[328]; 
    assign layer_0[6037] = in[437] ^ in[512]; 
    assign layer_0[6038] = in[763]; 
    assign layer_0[6039] = in[610] | in[88]; 
    assign layer_0[6040] = ~in[756]; 
    assign layer_0[6041] = in[401] & in[341]; 
    assign layer_0[6042] = in[466] ^ in[375]; 
    assign layer_0[6043] = ~in[585]; 
    assign layer_0[6044] = ~(in[205] | in[467]); 
    assign layer_0[6045] = ~in[150] | (in[150] & in[190]); 
    assign layer_0[6046] = in[261] ^ in[618]; 
    assign layer_0[6047] = in[50] ^ in[632]; 
    assign layer_0[6048] = ~in[619]; 
    assign layer_0[6049] = 1'b1; 
    assign layer_0[6050] = ~(in[95] | in[663]); 
    assign layer_0[6051] = ~(in[587] ^ in[634]); 
    assign layer_0[6052] = 1'b1; 
    assign layer_0[6053] = in[602] | in[508]; 
    assign layer_0[6054] = in[651] | in[583]; 
    assign layer_0[6055] = in[445] | in[608]; 
    assign layer_0[6056] = ~(in[743] ^ in[339]); 
    assign layer_0[6057] = ~in[61] | (in[420] & in[61]); 
    assign layer_0[6058] = in[664] & in[615]; 
    assign layer_0[6059] = in[76]; 
    assign layer_0[6060] = ~(in[19] ^ in[313]); 
    assign layer_0[6061] = ~in[372] | (in[372] & in[739]); 
    assign layer_0[6062] = ~in[81] | (in[81] & in[679]); 
    assign layer_0[6063] = ~(in[69] ^ in[671]); 
    assign layer_0[6064] = in[494] | in[307]; 
    assign layer_0[6065] = in[187] & ~in[579]; 
    assign layer_0[6066] = ~(in[388] ^ in[474]); 
    assign layer_0[6067] = in[222]; 
    assign layer_0[6068] = ~in[66]; 
    assign layer_0[6069] = ~(in[599] ^ in[759]); 
    assign layer_0[6070] = in[634]; 
    assign layer_0[6071] = in[308]; 
    assign layer_0[6072] = in[258] | in[534]; 
    assign layer_0[6073] = ~(in[685] ^ in[492]); 
    assign layer_0[6074] = in[427]; 
    assign layer_0[6075] = in[108] ^ in[195]; 
    assign layer_0[6076] = ~in[29] | (in[29] & in[668]); 
    assign layer_0[6077] = in[667]; 
    assign layer_0[6078] = in[83] | in[309]; 
    assign layer_0[6079] = in[445] & ~in[322]; 
    assign layer_0[6080] = in[40] & in[475]; 
    assign layer_0[6081] = in[409] & ~in[652]; 
    assign layer_0[6082] = in[62] & ~in[722]; 
    assign layer_0[6083] = ~(in[262] | in[317]); 
    assign layer_0[6084] = ~in[449]; 
    assign layer_0[6085] = ~(in[330] ^ in[501]); 
    assign layer_0[6086] = ~in[124]; 
    assign layer_0[6087] = ~in[712] | (in[712] & in[413]); 
    assign layer_0[6088] = ~in[604] | (in[604] & in[590]); 
    assign layer_0[6089] = in[641]; 
    assign layer_0[6090] = ~(in[64] ^ in[311]); 
    assign layer_0[6091] = in[104] ^ in[114]; 
    assign layer_0[6092] = ~in[500] | (in[500] & in[670]); 
    assign layer_0[6093] = ~in[554] | (in[34] & in[554]); 
    assign layer_0[6094] = in[717] & in[714]; 
    assign layer_0[6095] = ~in[246] | (in[583] & in[246]); 
    assign layer_0[6096] = ~(in[536] & in[428]); 
    assign layer_0[6097] = in[641] ^ in[314]; 
    assign layer_0[6098] = in[535] ^ in[531]; 
    assign layer_0[6099] = ~(in[653] & in[43]); 
    assign layer_0[6100] = in[81]; 
    assign layer_0[6101] = ~in[583] | (in[538] & in[583]); 
    assign layer_0[6102] = ~(in[538] ^ in[355]); 
    assign layer_0[6103] = ~(in[651] ^ in[45]); 
    assign layer_0[6104] = ~(in[709] ^ in[629]); 
    assign layer_0[6105] = ~in[712] | (in[19] & in[712]); 
    assign layer_0[6106] = in[583] & ~in[406]; 
    assign layer_0[6107] = ~in[310] | (in[309] & in[310]); 
    assign layer_0[6108] = ~(in[623] | in[728]); 
    assign layer_0[6109] = in[363] & in[438]; 
    assign layer_0[6110] = ~in[457]; 
    assign layer_0[6111] = ~(in[744] ^ in[692]); 
    assign layer_0[6112] = in[476] ^ in[597]; 
    assign layer_0[6113] = in[60] ^ in[9]; 
    assign layer_0[6114] = ~in[696]; 
    assign layer_0[6115] = ~(in[221] ^ in[355]); 
    assign layer_0[6116] = ~(in[222] & in[683]); 
    assign layer_0[6117] = ~(in[70] ^ in[97]); 
    assign layer_0[6118] = ~in[519]; 
    assign layer_0[6119] = ~(in[506] | in[644]); 
    assign layer_0[6120] = ~(in[3] ^ in[632]); 
    assign layer_0[6121] = in[339] ^ in[261]; 
    assign layer_0[6122] = in[282] & ~in[263]; 
    assign layer_0[6123] = in[454] & ~in[255]; 
    assign layer_0[6124] = in[474] | in[443]; 
    assign layer_0[6125] = in[641] & ~in[693]; 
    assign layer_0[6126] = in[202] & in[149]; 
    assign layer_0[6127] = in[614] & ~in[411]; 
    assign layer_0[6128] = ~(in[223] | in[112]); 
    assign layer_0[6129] = ~in[641]; 
    assign layer_0[6130] = ~in[300] | (in[677] & in[300]); 
    assign layer_0[6131] = ~(in[682] ^ in[680]); 
    assign layer_0[6132] = ~(in[253] ^ in[660]); 
    assign layer_0[6133] = in[376] & in[598]; 
    assign layer_0[6134] = ~in[397] | (in[397] & in[143]); 
    assign layer_0[6135] = ~in[125] | (in[209] & in[125]); 
    assign layer_0[6136] = in[663] & ~in[522]; 
    assign layer_0[6137] = ~in[693] | (in[419] & in[693]); 
    assign layer_0[6138] = ~in[472] | (in[10] & in[472]); 
    assign layer_0[6139] = ~(in[33] & in[355]); 
    assign layer_0[6140] = 1'b1; 
    assign layer_0[6141] = ~(in[254] & in[579]); 
    assign layer_0[6142] = in[534] | in[34]; 
    assign layer_0[6143] = in[716] & ~in[645]; 
    assign layer_0[6144] = ~(in[175] | in[75]); 
    assign layer_0[6145] = ~in[475] | (in[533] & in[475]); 
    assign layer_0[6146] = ~in[550] | (in[550] & in[623]); 
    assign layer_0[6147] = in[262] ^ in[568]; 
    assign layer_0[6148] = in[759] ^ in[711]; 
    assign layer_0[6149] = ~(in[767] ^ in[52]); 
    assign layer_0[6150] = in[246]; 
    assign layer_0[6151] = ~(in[674] ^ in[452]); 
    assign layer_0[6152] = ~(in[729] ^ in[237]); 
    assign layer_0[6153] = ~(in[606] ^ in[63]); 
    assign layer_0[6154] = ~(in[215] ^ in[476]); 
    assign layer_0[6155] = in[360]; 
    assign layer_0[6156] = in[62] ^ in[613]; 
    assign layer_0[6157] = ~(in[448] ^ in[614]); 
    assign layer_0[6158] = ~(in[636] ^ in[300]); 
    assign layer_0[6159] = in[314] | in[748]; 
    assign layer_0[6160] = ~in[95]; 
    assign layer_0[6161] = in[733] | in[241]; 
    assign layer_0[6162] = ~(in[565] | in[260]); 
    assign layer_0[6163] = in[501] ^ in[107]; 
    assign layer_0[6164] = in[314] ^ in[619]; 
    assign layer_0[6165] = ~(in[459] | in[723]); 
    assign layer_0[6166] = ~(in[709] & in[222]); 
    assign layer_0[6167] = ~(in[435] & in[252]); 
    assign layer_0[6168] = in[619] & ~in[658]; 
    assign layer_0[6169] = in[514] ^ in[563]; 
    assign layer_0[6170] = ~(in[268] ^ in[60]); 
    assign layer_0[6171] = in[535]; 
    assign layer_0[6172] = in[692]; 
    assign layer_0[6173] = in[388] & in[446]; 
    assign layer_0[6174] = in[714] ^ in[227]; 
    assign layer_0[6175] = ~(in[171] ^ in[582]); 
    assign layer_0[6176] = ~(in[381] & in[345]); 
    assign layer_0[6177] = in[261]; 
    assign layer_0[6178] = ~in[633]; 
    assign layer_0[6179] = in[356] & ~in[504]; 
    assign layer_0[6180] = ~(in[650] ^ in[266]); 
    assign layer_0[6181] = ~(in[488] | in[204]); 
    assign layer_0[6182] = ~(in[96] ^ in[317]); 
    assign layer_0[6183] = ~(in[475] ^ in[435]); 
    assign layer_0[6184] = ~(in[698] ^ in[629]); 
    assign layer_0[6185] = ~(in[349] | in[270]); 
    assign layer_0[6186] = ~(in[267] ^ in[156]); 
    assign layer_0[6187] = in[483]; 
    assign layer_0[6188] = ~in[419] | (in[478] & in[419]); 
    assign layer_0[6189] = ~in[445] | (in[445] & in[655]); 
    assign layer_0[6190] = ~in[636]; 
    assign layer_0[6191] = ~in[628] | (in[183] & in[628]); 
    assign layer_0[6192] = in[408] ^ in[54]; 
    assign layer_0[6193] = ~(in[519] ^ in[315]); 
    assign layer_0[6194] = in[686] & ~in[361]; 
    assign layer_0[6195] = ~in[317]; 
    assign layer_0[6196] = in[729]; 
    assign layer_0[6197] = in[127] & ~in[341]; 
    assign layer_0[6198] = in[414] ^ in[215]; 
    assign layer_0[6199] = ~in[77]; 
    assign layer_0[6200] = in[221] & in[96]; 
    assign layer_0[6201] = ~(in[683] | in[600]); 
    assign layer_0[6202] = ~in[39]; 
    assign layer_0[6203] = ~(in[468] ^ in[34]); 
    assign layer_0[6204] = ~(in[699] ^ in[484]); 
    assign layer_0[6205] = ~in[75] | (in[75] & in[463]); 
    assign layer_0[6206] = in[322]; 
    assign layer_0[6207] = in[347]; 
    assign layer_0[6208] = ~(in[192] | in[450]); 
    assign layer_0[6209] = ~(in[668] ^ in[729]); 
    assign layer_0[6210] = ~in[288]; 
    assign layer_0[6211] = ~(in[122] & in[151]); 
    assign layer_0[6212] = ~in[391] | (in[391] & in[398]); 
    assign layer_0[6213] = ~(in[594] | in[596]); 
    assign layer_0[6214] = ~(in[242] & in[114]); 
    assign layer_0[6215] = in[657] ^ in[55]; 
    assign layer_0[6216] = in[351] & ~in[734]; 
    assign layer_0[6217] = ~in[65]; 
    assign layer_0[6218] = in[728]; 
    assign layer_0[6219] = ~in[145] | (in[86] & in[145]); 
    assign layer_0[6220] = ~(in[611] | in[550]); 
    assign layer_0[6221] = in[177]; 
    assign layer_0[6222] = ~(in[729] & in[300]); 
    assign layer_0[6223] = ~(in[467] ^ in[160]); 
    assign layer_0[6224] = ~(in[641] ^ in[648]); 
    assign layer_0[6225] = in[307] & ~in[682]; 
    assign layer_0[6226] = ~in[759]; 
    assign layer_0[6227] = ~in[242] | (in[644] & in[242]); 
    assign layer_0[6228] = ~(in[62] ^ in[643]); 
    assign layer_0[6229] = ~in[420]; 
    assign layer_0[6230] = ~in[346] | (in[129] & in[346]); 
    assign layer_0[6231] = in[345] | in[618]; 
    assign layer_0[6232] = in[242] ^ in[98]; 
    assign layer_0[6233] = ~in[11]; 
    assign layer_0[6234] = ~(in[644] ^ in[243]); 
    assign layer_0[6235] = in[647] ^ in[633]; 
    assign layer_0[6236] = in[65] & ~in[702]; 
    assign layer_0[6237] = ~(in[354] | in[555]); 
    assign layer_0[6238] = 1'b1; 
    assign layer_0[6239] = in[615] | in[508]; 
    assign layer_0[6240] = ~(in[535] ^ in[563]); 
    assign layer_0[6241] = ~(in[187] & in[247]); 
    assign layer_0[6242] = in[694] & ~in[159]; 
    assign layer_0[6243] = ~(in[192] | in[654]); 
    assign layer_0[6244] = in[387] & in[77]; 
    assign layer_0[6245] = in[276] ^ in[10]; 
    assign layer_0[6246] = in[373] ^ in[202]; 
    assign layer_0[6247] = ~(in[57] ^ in[646]); 
    assign layer_0[6248] = ~(in[66] ^ in[293]); 
    assign layer_0[6249] = in[240] ^ in[248]; 
    assign layer_0[6250] = in[308] & ~in[28]; 
    assign layer_0[6251] = in[698] ^ in[331]; 
    assign layer_0[6252] = ~(in[597] ^ in[693]); 
    assign layer_0[6253] = ~(in[636] ^ in[665]); 
    assign layer_0[6254] = ~(in[468] ^ in[602]); 
    assign layer_0[6255] = in[1] & ~in[125]; 
    assign layer_0[6256] = ~in[717]; 
    assign layer_0[6257] = ~in[210]; 
    assign layer_0[6258] = in[712] & ~in[253]; 
    assign layer_0[6259] = ~(in[594] & in[7]); 
    assign layer_0[6260] = in[99] & ~in[574]; 
    assign layer_0[6261] = ~(in[121] & in[655]); 
    assign layer_0[6262] = ~in[291] | (in[291] & in[274]); 
    assign layer_0[6263] = ~(in[538] ^ in[439]); 
    assign layer_0[6264] = in[615] & ~in[671]; 
    assign layer_0[6265] = in[296] ^ in[19]; 
    assign layer_0[6266] = in[419] & ~in[242]; 
    assign layer_0[6267] = in[399] ^ in[267]; 
    assign layer_0[6268] = ~in[51]; 
    assign layer_0[6269] = in[412] | in[692]; 
    assign layer_0[6270] = ~(in[442] ^ in[753]); 
    assign layer_0[6271] = in[289]; 
    assign layer_0[6272] = in[474] ^ in[477]; 
    assign layer_0[6273] = ~(in[491] ^ in[549]); 
    assign layer_0[6274] = ~(in[743] | in[475]); 
    assign layer_0[6275] = in[684] ^ in[371]; 
    assign layer_0[6276] = in[251] ^ in[521]; 
    assign layer_0[6277] = in[277] & in[597]; 
    assign layer_0[6278] = in[66] | in[570]; 
    assign layer_0[6279] = ~(in[664] ^ in[504]); 
    assign layer_0[6280] = in[692] ^ in[661]; 
    assign layer_0[6281] = ~(in[503] | in[29]); 
    assign layer_0[6282] = ~in[201] | (in[194] & in[201]); 
    assign layer_0[6283] = ~(in[586] ^ in[340]); 
    assign layer_0[6284] = in[459] ^ in[569]; 
    assign layer_0[6285] = ~(in[23] ^ in[446]); 
    assign layer_0[6286] = ~(in[320] | in[154]); 
    assign layer_0[6287] = ~in[727] | (in[727] & in[597]); 
    assign layer_0[6288] = in[440]; 
    assign layer_0[6289] = ~(in[344] ^ in[119]); 
    assign layer_0[6290] = ~in[537]; 
    assign layer_0[6291] = in[238] | in[416]; 
    assign layer_0[6292] = in[671] | in[494]; 
    assign layer_0[6293] = ~in[206] | (in[672] & in[206]); 
    assign layer_0[6294] = in[163] ^ in[454]; 
    assign layer_0[6295] = ~in[163]; 
    assign layer_0[6296] = in[101] ^ in[311]; 
    assign layer_0[6297] = ~in[470] | (in[257] & in[470]); 
    assign layer_0[6298] = ~(in[331] ^ in[266]); 
    assign layer_0[6299] = ~in[590]; 
    assign layer_0[6300] = in[316] ^ in[683]; 
    assign layer_0[6301] = in[22] ^ in[238]; 
    assign layer_0[6302] = in[192] ^ in[358]; 
    assign layer_0[6303] = ~in[386] | (in[386] & in[684]); 
    assign layer_0[6304] = ~(in[513] | in[199]); 
    assign layer_0[6305] = in[110]; 
    assign layer_0[6306] = in[393] & ~in[566]; 
    assign layer_0[6307] = ~in[193]; 
    assign layer_0[6308] = in[572] | in[580]; 
    assign layer_0[6309] = ~(in[569] ^ in[570]); 
    assign layer_0[6310] = ~(in[300] ^ in[615]); 
    assign layer_0[6311] = in[695] & in[411]; 
    assign layer_0[6312] = in[599] | in[160]; 
    assign layer_0[6313] = in[437] | in[8]; 
    assign layer_0[6314] = in[612] ^ in[613]; 
    assign layer_0[6315] = ~(in[633] ^ in[665]); 
    assign layer_0[6316] = ~in[356]; 
    assign layer_0[6317] = in[519] & ~in[18]; 
    assign layer_0[6318] = ~(in[351] ^ in[516]); 
    assign layer_0[6319] = in[536] ^ in[551]; 
    assign layer_0[6320] = in[588] ^ in[567]; 
    assign layer_0[6321] = ~in[101]; 
    assign layer_0[6322] = ~in[623]; 
    assign layer_0[6323] = ~(in[252] ^ in[428]); 
    assign layer_0[6324] = ~in[614] | (in[635] & in[614]); 
    assign layer_0[6325] = in[489] | in[716]; 
    assign layer_0[6326] = in[283] & ~in[275]; 
    assign layer_0[6327] = ~(in[248] ^ in[659]); 
    assign layer_0[6328] = ~(in[194] ^ in[98]); 
    assign layer_0[6329] = ~(in[409] ^ in[424]); 
    assign layer_0[6330] = in[19] & in[423]; 
    assign layer_0[6331] = in[46] & in[94]; 
    assign layer_0[6332] = in[266] | in[13]; 
    assign layer_0[6333] = ~(in[399] | in[627]); 
    assign layer_0[6334] = in[681] ^ in[170]; 
    assign layer_0[6335] = in[301] ^ in[6]; 
    assign layer_0[6336] = in[390] & in[588]; 
    assign layer_0[6337] = in[51] & ~in[46]; 
    assign layer_0[6338] = in[274] | in[709]; 
    assign layer_0[6339] = ~(in[629] | in[629]); 
    assign layer_0[6340] = in[656] & ~in[97]; 
    assign layer_0[6341] = in[325]; 
    assign layer_0[6342] = ~(in[26] ^ in[616]); 
    assign layer_0[6343] = in[264] ^ in[618]; 
    assign layer_0[6344] = ~in[679] | (in[679] & in[602]); 
    assign layer_0[6345] = in[159] ^ in[745]; 
    assign layer_0[6346] = ~(in[583] ^ in[726]); 
    assign layer_0[6347] = in[118] & in[698]; 
    assign layer_0[6348] = in[407] & in[205]; 
    assign layer_0[6349] = in[669] ^ in[507]; 
    assign layer_0[6350] = in[138] ^ in[80]; 
    assign layer_0[6351] = in[53] & ~in[501]; 
    assign layer_0[6352] = in[221] & ~in[17]; 
    assign layer_0[6353] = in[342] & ~in[521]; 
    assign layer_0[6354] = in[111] | in[265]; 
    assign layer_0[6355] = in[236] ^ in[724]; 
    assign layer_0[6356] = ~in[418]; 
    assign layer_0[6357] = in[293]; 
    assign layer_0[6358] = in[690] & in[209]; 
    assign layer_0[6359] = in[276]; 
    assign layer_0[6360] = ~(in[491] ^ in[238]); 
    assign layer_0[6361] = ~(in[505] & in[648]); 
    assign layer_0[6362] = in[84]; 
    assign layer_0[6363] = ~(in[199] ^ in[314]); 
    assign layer_0[6364] = ~in[680] | (in[680] & in[226]); 
    assign layer_0[6365] = ~(in[402] ^ in[158]); 
    assign layer_0[6366] = in[76] & ~in[465]; 
    assign layer_0[6367] = in[614] ^ in[483]; 
    assign layer_0[6368] = 1'b0; 
    assign layer_0[6369] = ~(in[314] | in[554]); 
    assign layer_0[6370] = in[633] & in[617]; 
    assign layer_0[6371] = in[617] ^ in[652]; 
    assign layer_0[6372] = ~(in[194] ^ in[372]); 
    assign layer_0[6373] = ~in[351] | (in[351] & in[565]); 
    assign layer_0[6374] = ~in[596]; 
    assign layer_0[6375] = ~(in[636] ^ in[746]); 
    assign layer_0[6376] = in[253] ^ in[34]; 
    assign layer_0[6377] = in[726] ^ in[364]; 
    assign layer_0[6378] = in[102] & ~in[322]; 
    assign layer_0[6379] = in[149] & in[262]; 
    assign layer_0[6380] = ~in[49]; 
    assign layer_0[6381] = in[19] ^ in[677]; 
    assign layer_0[6382] = in[177] | in[353]; 
    assign layer_0[6383] = in[318] ^ in[659]; 
    assign layer_0[6384] = in[67] & in[451]; 
    assign layer_0[6385] = ~(in[353] ^ in[720]); 
    assign layer_0[6386] = in[268] ^ in[463]; 
    assign layer_0[6387] = in[44] ^ in[308]; 
    assign layer_0[6388] = in[490] & in[292]; 
    assign layer_0[6389] = ~(in[758] ^ in[193]); 
    assign layer_0[6390] = in[664] & ~in[277]; 
    assign layer_0[6391] = ~(in[712] | in[611]); 
    assign layer_0[6392] = ~in[642] | (in[479] & in[642]); 
    assign layer_0[6393] = ~in[581] | (in[581] & in[730]); 
    assign layer_0[6394] = ~(in[58] & in[755]); 
    assign layer_0[6395] = ~in[357] | (in[381] & in[357]); 
    assign layer_0[6396] = ~in[587]; 
    assign layer_0[6397] = in[667] ^ in[665]; 
    assign layer_0[6398] = ~in[468]; 
    assign layer_0[6399] = ~in[352] | (in[352] & in[332]); 
    assign layer_0[6400] = ~in[135] | (in[347] & in[135]); 
    assign layer_0[6401] = ~in[682] | (in[583] & in[682]); 
    assign layer_0[6402] = ~in[202] | (in[544] & in[202]); 
    assign layer_0[6403] = in[583] ^ in[292]; 
    assign layer_0[6404] = ~(in[613] | in[703]); 
    assign layer_0[6405] = in[619] ^ in[730]; 
    assign layer_0[6406] = in[254] ^ in[221]; 
    assign layer_0[6407] = ~in[659]; 
    assign layer_0[6408] = in[437] & ~in[450]; 
    assign layer_0[6409] = in[82] & ~in[98]; 
    assign layer_0[6410] = ~in[195]; 
    assign layer_0[6411] = in[324] & ~in[518]; 
    assign layer_0[6412] = in[656] ^ in[669]; 
    assign layer_0[6413] = in[138] & in[388]; 
    assign layer_0[6414] = ~in[471]; 
    assign layer_0[6415] = ~in[184] | (in[327] & in[184]); 
    assign layer_0[6416] = ~(in[65] ^ in[259]); 
    assign layer_0[6417] = ~(in[685] ^ in[134]); 
    assign layer_0[6418] = ~(in[681] | in[603]); 
    assign layer_0[6419] = ~(in[629] | in[635]); 
    assign layer_0[6420] = in[340]; 
    assign layer_0[6421] = ~in[279]; 
    assign layer_0[6422] = in[373] ^ in[716]; 
    assign layer_0[6423] = in[227] ^ in[403]; 
    assign layer_0[6424] = ~in[23] | (in[240] & in[23]); 
    assign layer_0[6425] = ~(in[1] ^ in[632]); 
    assign layer_0[6426] = ~in[98]; 
    assign layer_0[6427] = ~(in[296] ^ in[129]); 
    assign layer_0[6428] = in[685] ^ in[572]; 
    assign layer_0[6429] = ~in[340] | (in[614] & in[340]); 
    assign layer_0[6430] = ~(in[299] ^ in[733]); 
    assign layer_0[6431] = in[425] ^ in[743]; 
    assign layer_0[6432] = ~(in[157] ^ in[631]); 
    assign layer_0[6433] = ~(in[596] | in[197]); 
    assign layer_0[6434] = in[60] ^ in[622]; 
    assign layer_0[6435] = ~in[684] | (in[630] & in[684]); 
    assign layer_0[6436] = in[49] | in[562]; 
    assign layer_0[6437] = ~in[392] | (in[514] & in[392]); 
    assign layer_0[6438] = ~in[700]; 
    assign layer_0[6439] = ~(in[141] & in[5]); 
    assign layer_0[6440] = ~(in[628] ^ in[316]); 
    assign layer_0[6441] = ~(in[476] ^ in[264]); 
    assign layer_0[6442] = ~in[732] | (in[691] & in[732]); 
    assign layer_0[6443] = 1'b1; 
    assign layer_0[6444] = in[726] | in[266]; 
    assign layer_0[6445] = in[210]; 
    assign layer_0[6446] = ~(in[83] ^ in[673]); 
    assign layer_0[6447] = ~in[261]; 
    assign layer_0[6448] = in[639] | in[748]; 
    assign layer_0[6449] = in[145] ^ in[111]; 
    assign layer_0[6450] = in[666] ^ in[452]; 
    assign layer_0[6451] = in[410] ^ in[555]; 
    assign layer_0[6452] = in[236] & ~in[347]; 
    assign layer_0[6453] = ~(in[110] ^ in[651]); 
    assign layer_0[6454] = ~in[194] | (in[703] & in[194]); 
    assign layer_0[6455] = in[94] & in[160]; 
    assign layer_0[6456] = ~in[243]; 
    assign layer_0[6457] = in[370] | in[535]; 
    assign layer_0[6458] = in[279] | in[352]; 
    assign layer_0[6459] = ~in[659]; 
    assign layer_0[6460] = in[581]; 
    assign layer_0[6461] = ~in[501] | (in[501] & in[625]); 
    assign layer_0[6462] = ~in[279] | (in[279] & in[262]); 
    assign layer_0[6463] = ~in[643] | (in[643] & in[505]); 
    assign layer_0[6464] = in[671] ^ in[614]; 
    assign layer_0[6465] = ~(in[565] | in[271]); 
    assign layer_0[6466] = in[87] & in[25]; 
    assign layer_0[6467] = ~(in[314] | in[630]); 
    assign layer_0[6468] = ~(in[244] | in[160]); 
    assign layer_0[6469] = in[747] ^ in[682]; 
    assign layer_0[6470] = in[712] ^ in[162]; 
    assign layer_0[6471] = in[167] | in[183]; 
    assign layer_0[6472] = in[223] ^ in[255]; 
    assign layer_0[6473] = ~(in[74] & in[80]); 
    assign layer_0[6474] = in[327] & in[13]; 
    assign layer_0[6475] = in[435]; 
    assign layer_0[6476] = ~in[11]; 
    assign layer_0[6477] = in[627] & ~in[501]; 
    assign layer_0[6478] = ~in[434]; 
    assign layer_0[6479] = in[55] ^ in[384]; 
    assign layer_0[6480] = ~in[56] | (in[56] & in[599]); 
    assign layer_0[6481] = in[310] & ~in[49]; 
    assign layer_0[6482] = ~(in[335] | in[669]); 
    assign layer_0[6483] = ~(in[569] | in[282]); 
    assign layer_0[6484] = ~in[11] | (in[287] & in[11]); 
    assign layer_0[6485] = ~(in[158] ^ in[746]); 
    assign layer_0[6486] = in[708]; 
    assign layer_0[6487] = ~(in[51] ^ in[272]); 
    assign layer_0[6488] = in[520] ^ in[396]; 
    assign layer_0[6489] = in[714] ^ in[518]; 
    assign layer_0[6490] = in[471]; 
    assign layer_0[6491] = in[541] ^ in[230]; 
    assign layer_0[6492] = ~(in[222] | in[349]); 
    assign layer_0[6493] = ~(in[574] | in[160]); 
    assign layer_0[6494] = ~(in[52] & in[620]); 
    assign layer_0[6495] = in[34] | in[445]; 
    assign layer_0[6496] = in[329] & ~in[554]; 
    assign layer_0[6497] = in[34] | in[242]; 
    assign layer_0[6498] = in[471] | in[59]; 
    assign layer_0[6499] = ~in[306] | (in[306] & in[81]); 
    assign layer_0[6500] = 1'b0; 
    assign layer_0[6501] = ~in[69]; 
    assign layer_0[6502] = in[663] & ~in[632]; 
    assign layer_0[6503] = in[695] ^ in[710]; 
    assign layer_0[6504] = ~(in[336] | in[124]); 
    assign layer_0[6505] = in[614] ^ in[338]; 
    assign layer_0[6506] = ~in[553]; 
    assign layer_0[6507] = in[180] & ~in[509]; 
    assign layer_0[6508] = in[22] & ~in[143]; 
    assign layer_0[6509] = in[370] ^ in[46]; 
    assign layer_0[6510] = in[628] & in[237]; 
    assign layer_0[6511] = ~in[9] | (in[9] & in[227]); 
    assign layer_0[6512] = in[112] & in[21]; 
    assign layer_0[6513] = ~in[331] | (in[622] & in[331]); 
    assign layer_0[6514] = ~in[740]; 
    assign layer_0[6515] = in[711] & ~in[411]; 
    assign layer_0[6516] = in[80] ^ in[50]; 
    assign layer_0[6517] = ~in[150] | (in[150] & in[611]); 
    assign layer_0[6518] = ~(in[452] ^ in[475]); 
    assign layer_0[6519] = ~(in[439] | in[17]); 
    assign layer_0[6520] = in[445]; 
    assign layer_0[6521] = in[640] | in[325]; 
    assign layer_0[6522] = ~(in[192] | in[358]); 
    assign layer_0[6523] = ~(in[70] ^ in[197]); 
    assign layer_0[6524] = in[281] & ~in[264]; 
    assign layer_0[6525] = in[662] | in[198]; 
    assign layer_0[6526] = in[586]; 
    assign layer_0[6527] = ~(in[43] & in[433]); 
    assign layer_0[6528] = ~(in[610] & in[200]); 
    assign layer_0[6529] = ~(in[143] ^ in[606]); 
    assign layer_0[6530] = ~(in[606] | in[30]); 
    assign layer_0[6531] = in[648] ^ in[43]; 
    assign layer_0[6532] = ~(in[64] | in[667]); 
    assign layer_0[6533] = ~(in[679] ^ in[86]); 
    assign layer_0[6534] = in[646] & ~in[739]; 
    assign layer_0[6535] = ~in[359] | (in[299] & in[359]); 
    assign layer_0[6536] = in[552] & ~in[757]; 
    assign layer_0[6537] = in[337]; 
    assign layer_0[6538] = in[403]; 
    assign layer_0[6539] = in[170] & in[385]; 
    assign layer_0[6540] = in[584] & ~in[660]; 
    assign layer_0[6541] = in[11] ^ in[316]; 
    assign layer_0[6542] = ~in[464] | (in[353] & in[464]); 
    assign layer_0[6543] = ~(in[432] ^ in[201]); 
    assign layer_0[6544] = ~(in[638] ^ in[676]); 
    assign layer_0[6545] = ~in[696]; 
    assign layer_0[6546] = in[265]; 
    assign layer_0[6547] = ~in[161] | (in[275] & in[161]); 
    assign layer_0[6548] = in[611] & in[260]; 
    assign layer_0[6549] = ~in[223]; 
    assign layer_0[6550] = in[409] & in[563]; 
    assign layer_0[6551] = ~(in[380] ^ in[376]); 
    assign layer_0[6552] = 1'b1; 
    assign layer_0[6553] = in[225] | in[581]; 
    assign layer_0[6554] = in[423] & ~in[401]; 
    assign layer_0[6555] = ~in[476] | (in[386] & in[476]); 
    assign layer_0[6556] = ~(in[373] ^ in[729]); 
    assign layer_0[6557] = in[307]; 
    assign layer_0[6558] = 1'b0; 
    assign layer_0[6559] = ~(in[422] ^ in[8]); 
    assign layer_0[6560] = in[117]; 
    assign layer_0[6561] = in[632] ^ in[267]; 
    assign layer_0[6562] = 1'b0; 
    assign layer_0[6563] = ~in[34]; 
    assign layer_0[6564] = in[122] & in[124]; 
    assign layer_0[6565] = ~in[366] | (in[366] & in[257]); 
    assign layer_0[6566] = ~(in[307] ^ in[651]); 
    assign layer_0[6567] = in[300] ^ in[265]; 
    assign layer_0[6568] = ~(in[354] ^ in[620]); 
    assign layer_0[6569] = ~(in[699] ^ in[586]); 
    assign layer_0[6570] = ~(in[644] ^ in[473]); 
    assign layer_0[6571] = ~(in[709] ^ in[694]); 
    assign layer_0[6572] = in[450] | in[161]; 
    assign layer_0[6573] = in[225] | in[757]; 
    assign layer_0[6574] = ~(in[404] ^ in[759]); 
    assign layer_0[6575] = in[323]; 
    assign layer_0[6576] = in[600] & ~in[28]; 
    assign layer_0[6577] = in[638] ^ in[689]; 
    assign layer_0[6578] = in[373] & ~in[682]; 
    assign layer_0[6579] = in[555] | in[570]; 
    assign layer_0[6580] = in[678] & ~in[692]; 
    assign layer_0[6581] = ~(in[234] & in[393]); 
    assign layer_0[6582] = ~(in[627] ^ in[619]); 
    assign layer_0[6583] = ~in[12] | (in[12] & in[62]); 
    assign layer_0[6584] = in[538] & ~in[472]; 
    assign layer_0[6585] = in[681]; 
    assign layer_0[6586] = in[299] ^ in[242]; 
    assign layer_0[6587] = in[681] ^ in[601]; 
    assign layer_0[6588] = in[296] | in[555]; 
    assign layer_0[6589] = ~(in[746] | in[301]); 
    assign layer_0[6590] = ~(in[491] ^ in[714]); 
    assign layer_0[6591] = in[350] & ~in[574]; 
    assign layer_0[6592] = in[654] ^ in[370]; 
    assign layer_0[6593] = ~in[34] | (in[34] & in[451]); 
    assign layer_0[6594] = in[459]; 
    assign layer_0[6595] = in[60] | in[655]; 
    assign layer_0[6596] = 1'b0; 
    assign layer_0[6597] = in[536] ^ in[533]; 
    assign layer_0[6598] = in[522]; 
    assign layer_0[6599] = ~(in[185] | in[56]); 
    assign layer_0[6600] = in[46] ^ in[36]; 
    assign layer_0[6601] = ~(in[635] ^ in[476]); 
    assign layer_0[6602] = in[21] & in[508]; 
    assign layer_0[6603] = ~in[389]; 
    assign layer_0[6604] = in[264] | in[609]; 
    assign layer_0[6605] = in[29] & in[131]; 
    assign layer_0[6606] = ~(in[214] ^ in[49]); 
    assign layer_0[6607] = ~(in[519] ^ in[484]); 
    assign layer_0[6608] = in[582] | in[696]; 
    assign layer_0[6609] = in[28] & ~in[472]; 
    assign layer_0[6610] = ~(in[693] ^ in[598]); 
    assign layer_0[6611] = ~(in[498] | in[550]); 
    assign layer_0[6612] = ~(in[662] ^ in[217]); 
    assign layer_0[6613] = in[522]; 
    assign layer_0[6614] = ~in[60] | (in[60] & in[9]); 
    assign layer_0[6615] = ~(in[740] ^ in[256]); 
    assign layer_0[6616] = in[194]; 
    assign layer_0[6617] = in[44] ^ in[436]; 
    assign layer_0[6618] = ~in[593]; 
    assign layer_0[6619] = in[711] & ~in[190]; 
    assign layer_0[6620] = ~(in[724] ^ in[485]); 
    assign layer_0[6621] = ~(in[567] ^ in[554]); 
    assign layer_0[6622] = ~(in[185] & in[354]); 
    assign layer_0[6623] = in[196] ^ in[508]; 
    assign layer_0[6624] = in[46]; 
    assign layer_0[6625] = in[268]; 
    assign layer_0[6626] = ~in[44] | (in[718] & in[44]); 
    assign layer_0[6627] = ~in[653] | (in[702] & in[653]); 
    assign layer_0[6628] = in[614] & ~in[696]; 
    assign layer_0[6629] = ~(in[542] & in[645]); 
    assign layer_0[6630] = in[124]; 
    assign layer_0[6631] = ~in[237] | (in[237] & in[260]); 
    assign layer_0[6632] = ~(in[278] | in[413]); 
    assign layer_0[6633] = ~(in[620] ^ in[694]); 
    assign layer_0[6634] = in[479] ^ in[378]; 
    assign layer_0[6635] = ~(in[484] ^ in[760]); 
    assign layer_0[6636] = in[77] & ~in[676]; 
    assign layer_0[6637] = ~(in[229] ^ in[597]); 
    assign layer_0[6638] = in[28] & ~in[548]; 
    assign layer_0[6639] = in[388] ^ in[175]; 
    assign layer_0[6640] = ~(in[665] ^ in[417]); 
    assign layer_0[6641] = in[715] ^ in[748]; 
    assign layer_0[6642] = ~in[216] | (in[216] & in[681]); 
    assign layer_0[6643] = in[310] ^ in[346]; 
    assign layer_0[6644] = in[328]; 
    assign layer_0[6645] = ~(in[113] ^ in[60]); 
    assign layer_0[6646] = in[603] | in[100]; 
    assign layer_0[6647] = ~(in[35] | in[158]); 
    assign layer_0[6648] = ~in[612] | (in[612] & in[717]); 
    assign layer_0[6649] = in[265]; 
    assign layer_0[6650] = ~in[379] | (in[379] & in[387]); 
    assign layer_0[6651] = ~(in[208] ^ in[187]); 
    assign layer_0[6652] = ~(in[494] | in[242]); 
    assign layer_0[6653] = in[476]; 
    assign layer_0[6654] = ~in[43]; 
    assign layer_0[6655] = in[10] | in[528]; 
    assign layer_0[6656] = in[707] & ~in[646]; 
    assign layer_0[6657] = ~(in[64] | in[700]); 
    assign layer_0[6658] = in[605] | in[283]; 
    assign layer_0[6659] = in[252] & ~in[293]; 
    assign layer_0[6660] = in[377] & ~in[304]; 
    assign layer_0[6661] = in[509] | in[277]; 
    assign layer_0[6662] = ~(in[158] & in[240]); 
    assign layer_0[6663] = in[100] & in[619]; 
    assign layer_0[6664] = in[631] & ~in[521]; 
    assign layer_0[6665] = ~in[298]; 
    assign layer_0[6666] = in[13] | in[342]; 
    assign layer_0[6667] = ~in[8]; 
    assign layer_0[6668] = ~(in[709] ^ in[675]); 
    assign layer_0[6669] = ~(in[470] ^ in[764]); 
    assign layer_0[6670] = in[265] & in[429]; 
    assign layer_0[6671] = in[15] & ~in[677]; 
    assign layer_0[6672] = in[698] ^ in[534]; 
    assign layer_0[6673] = ~(in[470] & in[465]); 
    assign layer_0[6674] = ~(in[284] & in[704]); 
    assign layer_0[6675] = in[78] & ~in[224]; 
    assign layer_0[6676] = in[492] ^ in[375]; 
    assign layer_0[6677] = in[280] & ~in[531]; 
    assign layer_0[6678] = ~(in[174] ^ in[340]); 
    assign layer_0[6679] = in[18] & ~in[573]; 
    assign layer_0[6680] = ~in[675]; 
    assign layer_0[6681] = in[700] & ~in[711]; 
    assign layer_0[6682] = ~in[672]; 
    assign layer_0[6683] = ~in[150] | (in[150] & in[498]); 
    assign layer_0[6684] = ~(in[301] ^ in[309]); 
    assign layer_0[6685] = 1'b1; 
    assign layer_0[6686] = ~(in[675] ^ in[498]); 
    assign layer_0[6687] = in[112]; 
    assign layer_0[6688] = in[221]; 
    assign layer_0[6689] = ~in[359]; 
    assign layer_0[6690] = ~(in[112] ^ in[56]); 
    assign layer_0[6691] = in[318] & ~in[438]; 
    assign layer_0[6692] = ~(in[572] | in[144]); 
    assign layer_0[6693] = in[714] ^ in[750]; 
    assign layer_0[6694] = in[420] & ~in[484]; 
    assign layer_0[6695] = ~(in[691] | in[198]); 
    assign layer_0[6696] = in[692]; 
    assign layer_0[6697] = in[17]; 
    assign layer_0[6698] = in[757] | in[264]; 
    assign layer_0[6699] = ~(in[134] | in[413]); 
    assign layer_0[6700] = in[628] | in[632]; 
    assign layer_0[6701] = in[533] ^ in[261]; 
    assign layer_0[6702] = in[552] ^ in[263]; 
    assign layer_0[6703] = ~(in[5] & in[409]); 
    assign layer_0[6704] = ~(in[347] ^ in[666]); 
    assign layer_0[6705] = in[429] ^ in[604]; 
    assign layer_0[6706] = ~(in[77] ^ in[594]); 
    assign layer_0[6707] = ~in[287] | (in[287] & in[347]); 
    assign layer_0[6708] = ~in[725] | (in[725] & in[301]); 
    assign layer_0[6709] = in[109] & in[643]; 
    assign layer_0[6710] = ~(in[45] | in[619]); 
    assign layer_0[6711] = ~(in[409] & in[436]); 
    assign layer_0[6712] = in[597] & in[254]; 
    assign layer_0[6713] = in[132] ^ in[230]; 
    assign layer_0[6714] = in[533] ^ in[208]; 
    assign layer_0[6715] = in[634]; 
    assign layer_0[6716] = ~in[43] | (in[710] & in[43]); 
    assign layer_0[6717] = in[488]; 
    assign layer_0[6718] = ~in[245] | (in[245] & in[619]); 
    assign layer_0[6719] = ~in[111] | (in[544] & in[111]); 
    assign layer_0[6720] = ~(in[396] | in[347]); 
    assign layer_0[6721] = ~(in[51] | in[528]); 
    assign layer_0[6722] = in[177] & ~in[65]; 
    assign layer_0[6723] = in[113] & ~in[318]; 
    assign layer_0[6724] = in[584] ^ in[337]; 
    assign layer_0[6725] = ~(in[280] & in[380]); 
    assign layer_0[6726] = ~(in[177] ^ in[429]); 
    assign layer_0[6727] = in[430]; 
    assign layer_0[6728] = ~in[8]; 
    assign layer_0[6729] = in[375] & ~in[611]; 
    assign layer_0[6730] = in[311] | in[461]; 
    assign layer_0[6731] = in[147] ^ in[409]; 
    assign layer_0[6732] = in[260]; 
    assign layer_0[6733] = in[63] & ~in[474]; 
    assign layer_0[6734] = ~(in[694] & in[82]); 
    assign layer_0[6735] = in[348] & in[628]; 
    assign layer_0[6736] = in[698] & ~in[293]; 
    assign layer_0[6737] = ~in[144] | (in[301] & in[144]); 
    assign layer_0[6738] = in[476] ^ in[189]; 
    assign layer_0[6739] = in[373] & in[611]; 
    assign layer_0[6740] = ~in[587] | (in[345] & in[587]); 
    assign layer_0[6741] = in[612]; 
    assign layer_0[6742] = ~in[602] | (in[533] & in[602]); 
    assign layer_0[6743] = in[264] & ~in[552]; 
    assign layer_0[6744] = ~in[466]; 
    assign layer_0[6745] = ~in[565] | (in[565] & in[490]); 
    assign layer_0[6746] = in[696]; 
    assign layer_0[6747] = in[264] & in[479]; 
    assign layer_0[6748] = ~in[605]; 
    assign layer_0[6749] = ~in[217] | (in[519] & in[217]); 
    assign layer_0[6750] = ~in[501] | (in[660] & in[501]); 
    assign layer_0[6751] = ~(in[296] & in[633]); 
    assign layer_0[6752] = in[724] | in[299]; 
    assign layer_0[6753] = ~in[8] | (in[8] & in[649]); 
    assign layer_0[6754] = in[475] ^ in[533]; 
    assign layer_0[6755] = in[207] & in[333]; 
    assign layer_0[6756] = ~(in[404] ^ in[746]); 
    assign layer_0[6757] = in[620]; 
    assign layer_0[6758] = in[476] | in[684]; 
    assign layer_0[6759] = ~(in[655] & in[671]); 
    assign layer_0[6760] = in[160] & ~in[383]; 
    assign layer_0[6761] = ~in[360]; 
    assign layer_0[6762] = ~(in[683] & in[602]); 
    assign layer_0[6763] = ~(in[645] ^ in[693]); 
    assign layer_0[6764] = ~(in[402] & in[48]); 
    assign layer_0[6765] = in[487] & ~in[318]; 
    assign layer_0[6766] = in[177] & in[328]; 
    assign layer_0[6767] = ~in[413]; 
    assign layer_0[6768] = ~(in[754] ^ in[10]); 
    assign layer_0[6769] = in[570] & ~in[733]; 
    assign layer_0[6770] = in[552] | in[746]; 
    assign layer_0[6771] = in[254] ^ in[678]; 
    assign layer_0[6772] = ~in[536] | (in[536] & in[621]); 
    assign layer_0[6773] = ~in[278]; 
    assign layer_0[6774] = ~in[521]; 
    assign layer_0[6775] = in[444] & in[8]; 
    assign layer_0[6776] = ~(in[312] | in[237]); 
    assign layer_0[6777] = ~(in[724] | in[97]); 
    assign layer_0[6778] = ~in[402]; 
    assign layer_0[6779] = ~in[162] | (in[162] & in[325]); 
    assign layer_0[6780] = in[77]; 
    assign layer_0[6781] = in[460] ^ in[157]; 
    assign layer_0[6782] = in[633] ^ in[300]; 
    assign layer_0[6783] = ~(in[470] ^ in[571]); 
    assign layer_0[6784] = in[76] & ~in[189]; 
    assign layer_0[6785] = ~in[377] | (in[377] & in[756]); 
    assign layer_0[6786] = in[28] | in[20]; 
    assign layer_0[6787] = in[65]; 
    assign layer_0[6788] = ~(in[633] | in[205]); 
    assign layer_0[6789] = in[508] ^ in[236]; 
    assign layer_0[6790] = in[484] ^ in[130]; 
    assign layer_0[6791] = in[458] ^ in[468]; 
    assign layer_0[6792] = in[242] | in[537]; 
    assign layer_0[6793] = in[266] ^ in[483]; 
    assign layer_0[6794] = in[715] ^ in[238]; 
    assign layer_0[6795] = in[604] ^ in[584]; 
    assign layer_0[6796] = ~in[650] | (in[46] & in[650]); 
    assign layer_0[6797] = in[356] & in[216]; 
    assign layer_0[6798] = in[331] & ~in[174]; 
    assign layer_0[6799] = in[750]; 
    assign layer_0[6800] = in[539] | in[174]; 
    assign layer_0[6801] = ~(in[305] ^ in[172]); 
    assign layer_0[6802] = ~(in[583] ^ in[586]); 
    assign layer_0[6803] = ~in[264] | (in[402] & in[264]); 
    assign layer_0[6804] = in[603] ^ in[697]; 
    assign layer_0[6805] = in[479] ^ in[603]; 
    assign layer_0[6806] = ~(in[146] & in[82]); 
    assign layer_0[6807] = in[622] | in[729]; 
    assign layer_0[6808] = ~(in[552] ^ in[253]); 
    assign layer_0[6809] = ~(in[360] ^ in[696]); 
    assign layer_0[6810] = in[677]; 
    assign layer_0[6811] = in[255] | in[589]; 
    assign layer_0[6812] = ~in[236] | (in[758] & in[236]); 
    assign layer_0[6813] = ~(in[15] ^ in[20]); 
    assign layer_0[6814] = ~in[434]; 
    assign layer_0[6815] = ~in[60] | (in[60] & in[566]); 
    assign layer_0[6816] = ~in[602] | (in[631] & in[602]); 
    assign layer_0[6817] = in[641] & ~in[693]; 
    assign layer_0[6818] = in[266]; 
    assign layer_0[6819] = ~(in[481] | in[529]); 
    assign layer_0[6820] = in[499] ^ in[628]; 
    assign layer_0[6821] = ~(in[393] | in[398]); 
    assign layer_0[6822] = in[190]; 
    assign layer_0[6823] = ~in[706]; 
    assign layer_0[6824] = in[95] & ~in[562]; 
    assign layer_0[6825] = in[158]; 
    assign layer_0[6826] = ~(in[207] & in[377]); 
    assign layer_0[6827] = ~(in[262] ^ in[81]); 
    assign layer_0[6828] = ~in[592]; 
    assign layer_0[6829] = ~(in[483] ^ in[486]); 
    assign layer_0[6830] = in[114] | in[209]; 
    assign layer_0[6831] = ~(in[371] & in[276]); 
    assign layer_0[6832] = ~in[689] | (in[689] & in[625]); 
    assign layer_0[6833] = ~(in[561] | in[143]); 
    assign layer_0[6834] = ~in[647] | (in[623] & in[647]); 
    assign layer_0[6835] = ~(in[10] ^ in[488]); 
    assign layer_0[6836] = ~in[250] | (in[250] & in[693]); 
    assign layer_0[6837] = in[477] | in[721]; 
    assign layer_0[6838] = in[504] & ~in[282]; 
    assign layer_0[6839] = ~in[728] | (in[42] & in[728]); 
    assign layer_0[6840] = in[164] & ~in[156]; 
    assign layer_0[6841] = in[219]; 
    assign layer_0[6842] = ~(in[708] ^ in[222]); 
    assign layer_0[6843] = in[675] & ~in[506]; 
    assign layer_0[6844] = ~(in[277] ^ in[395]); 
    assign layer_0[6845] = in[123] & ~in[99]; 
    assign layer_0[6846] = in[334]; 
    assign layer_0[6847] = ~in[132]; 
    assign layer_0[6848] = in[552] ^ in[588]; 
    assign layer_0[6849] = ~(in[718] | in[458]); 
    assign layer_0[6850] = ~(in[482] ^ in[332]); 
    assign layer_0[6851] = in[676] & in[177]; 
    assign layer_0[6852] = ~in[46]; 
    assign layer_0[6853] = ~in[210]; 
    assign layer_0[6854] = ~(in[632] ^ in[680]); 
    assign layer_0[6855] = ~in[459]; 
    assign layer_0[6856] = ~(in[614] ^ in[283]); 
    assign layer_0[6857] = ~(in[226] ^ in[457]); 
    assign layer_0[6858] = in[677]; 
    assign layer_0[6859] = in[146] & in[653]; 
    assign layer_0[6860] = in[698] & ~in[462]; 
    assign layer_0[6861] = in[729] ^ in[390]; 
    assign layer_0[6862] = in[184] & ~in[637]; 
    assign layer_0[6863] = ~in[571]; 
    assign layer_0[6864] = in[19] & in[436]; 
    assign layer_0[6865] = in[612] ^ in[301]; 
    assign layer_0[6866] = ~(in[760] ^ in[617]); 
    assign layer_0[6867] = 1'b0; 
    assign layer_0[6868] = in[730] | in[34]; 
    assign layer_0[6869] = in[276]; 
    assign layer_0[6870] = ~in[690]; 
    assign layer_0[6871] = ~(in[585] & in[598]); 
    assign layer_0[6872] = in[415] & ~in[693]; 
    assign layer_0[6873] = ~(in[356] & in[658]); 
    assign layer_0[6874] = in[746] ^ in[666]; 
    assign layer_0[6875] = ~in[253]; 
    assign layer_0[6876] = in[762] ^ in[598]; 
    assign layer_0[6877] = in[97] ^ in[644]; 
    assign layer_0[6878] = ~(in[245] & in[708]); 
    assign layer_0[6879] = in[57] | in[684]; 
    assign layer_0[6880] = in[343] & in[447]; 
    assign layer_0[6881] = in[252] & in[565]; 
    assign layer_0[6882] = in[457] ^ in[725]; 
    assign layer_0[6883] = ~(in[663] ^ in[661]); 
    assign layer_0[6884] = in[130] | in[563]; 
    assign layer_0[6885] = ~in[707]; 
    assign layer_0[6886] = in[174] & ~in[723]; 
    assign layer_0[6887] = ~(in[22] | in[509]); 
    assign layer_0[6888] = ~(in[627] & in[684]); 
    assign layer_0[6889] = ~(in[501] ^ in[12]); 
    assign layer_0[6890] = in[759] ^ in[645]; 
    assign layer_0[6891] = ~in[314]; 
    assign layer_0[6892] = in[486] ^ in[711]; 
    assign layer_0[6893] = in[473] & ~in[763]; 
    assign layer_0[6894] = in[426] & ~in[631]; 
    assign layer_0[6895] = ~(in[706] ^ in[4]); 
    assign layer_0[6896] = in[415] & ~in[291]; 
    assign layer_0[6897] = in[300] | in[638]; 
    assign layer_0[6898] = in[118]; 
    assign layer_0[6899] = in[3] ^ in[282]; 
    assign layer_0[6900] = ~(in[4] | in[461]); 
    assign layer_0[6901] = ~(in[678] ^ in[217]); 
    assign layer_0[6902] = ~in[324]; 
    assign layer_0[6903] = ~(in[368] | in[192]); 
    assign layer_0[6904] = ~(in[546] ^ in[300]); 
    assign layer_0[6905] = in[97] ^ in[668]; 
    assign layer_0[6906] = ~(in[276] | in[705]); 
    assign layer_0[6907] = in[600] | in[77]; 
    assign layer_0[6908] = in[728]; 
    assign layer_0[6909] = ~(in[507] ^ in[330]); 
    assign layer_0[6910] = ~in[51] | (in[564] & in[51]); 
    assign layer_0[6911] = in[334] | in[15]; 
    assign layer_0[6912] = ~(in[523] ^ in[301]); 
    assign layer_0[6913] = ~(in[662] | in[519]); 
    assign layer_0[6914] = in[359] & ~in[757]; 
    assign layer_0[6915] = in[355] ^ in[468]; 
    assign layer_0[6916] = ~(in[291] ^ in[81]); 
    assign layer_0[6917] = ~(in[442] | in[647]); 
    assign layer_0[6918] = ~in[582] | (in[411] & in[582]); 
    assign layer_0[6919] = ~(in[36] ^ in[692]); 
    assign layer_0[6920] = in[138] ^ in[343]; 
    assign layer_0[6921] = ~in[665]; 
    assign layer_0[6922] = in[323] & in[509]; 
    assign layer_0[6923] = ~in[162]; 
    assign layer_0[6924] = in[296] & ~in[466]; 
    assign layer_0[6925] = ~(in[742] ^ in[759]); 
    assign layer_0[6926] = ~(in[549] | in[357]); 
    assign layer_0[6927] = in[640] & ~in[275]; 
    assign layer_0[6928] = ~(in[518] ^ in[611]); 
    assign layer_0[6929] = ~(in[612] ^ in[261]); 
    assign layer_0[6930] = ~(in[556] ^ in[474]); 
    assign layer_0[6931] = in[222] ^ in[175]; 
    assign layer_0[6932] = ~in[159] | (in[159] & in[598]); 
    assign layer_0[6933] = in[53] | in[65]; 
    assign layer_0[6934] = ~(in[730] ^ in[727]); 
    assign layer_0[6935] = ~in[238]; 
    assign layer_0[6936] = in[19] ^ in[597]; 
    assign layer_0[6937] = ~in[499]; 
    assign layer_0[6938] = ~in[430]; 
    assign layer_0[6939] = ~(in[760] ^ in[761]); 
    assign layer_0[6940] = in[349]; 
    assign layer_0[6941] = ~in[458] | (in[232] & in[458]); 
    assign layer_0[6942] = in[232] & in[691]; 
    assign layer_0[6943] = ~in[483] | (in[483] & in[369]); 
    assign layer_0[6944] = ~(in[215] ^ in[384]); 
    assign layer_0[6945] = 1'b1; 
    assign layer_0[6946] = ~in[311] | (in[223] & in[311]); 
    assign layer_0[6947] = in[56] ^ in[334]; 
    assign layer_0[6948] = in[471] & ~in[662]; 
    assign layer_0[6949] = ~in[598]; 
    assign layer_0[6950] = ~(in[29] | in[296]); 
    assign layer_0[6951] = in[92] & ~in[690]; 
    assign layer_0[6952] = ~(in[740] ^ in[632]); 
    assign layer_0[6953] = in[509] | in[430]; 
    assign layer_0[6954] = ~(in[4] ^ in[460]); 
    assign layer_0[6955] = in[346] & ~in[271]; 
    assign layer_0[6956] = in[452] | in[601]; 
    assign layer_0[6957] = ~(in[422] & in[692]); 
    assign layer_0[6958] = ~in[633] | (in[235] & in[633]); 
    assign layer_0[6959] = ~(in[676] | in[355]); 
    assign layer_0[6960] = in[552] & ~in[45]; 
    assign layer_0[6961] = ~in[118] | (in[321] & in[118]); 
    assign layer_0[6962] = in[675] | in[614]; 
    assign layer_0[6963] = in[242] & ~in[357]; 
    assign layer_0[6964] = in[564] & in[587]; 
    assign layer_0[6965] = ~in[328] | (in[328] & in[335]); 
    assign layer_0[6966] = in[726] | in[259]; 
    assign layer_0[6967] = ~(in[36] ^ in[759]); 
    assign layer_0[6968] = in[302] | in[736]; 
    assign layer_0[6969] = ~in[231]; 
    assign layer_0[6970] = ~in[343] | (in[533] & in[343]); 
    assign layer_0[6971] = in[632] ^ in[630]; 
    assign layer_0[6972] = ~(in[250] & in[26]); 
    assign layer_0[6973] = ~in[245]; 
    assign layer_0[6974] = in[63]; 
    assign layer_0[6975] = ~in[563]; 
    assign layer_0[6976] = ~(in[191] ^ in[300]); 
    assign layer_0[6977] = in[551] ^ in[331]; 
    assign layer_0[6978] = in[198]; 
    assign layer_0[6979] = ~(in[595] ^ in[587]); 
    assign layer_0[6980] = ~(in[350] | in[754]); 
    assign layer_0[6981] = ~(in[655] | in[329]); 
    assign layer_0[6982] = in[162] | in[569]; 
    assign layer_0[6983] = ~(in[75] & in[326]); 
    assign layer_0[6984] = ~in[570]; 
    assign layer_0[6985] = in[383]; 
    assign layer_0[6986] = in[349] & in[611]; 
    assign layer_0[6987] = ~(in[724] ^ in[245]); 
    assign layer_0[6988] = in[433] & ~in[628]; 
    assign layer_0[6989] = in[177]; 
    assign layer_0[6990] = in[656] | in[45]; 
    assign layer_0[6991] = in[566] ^ in[568]; 
    assign layer_0[6992] = ~(in[631] ^ in[746]); 
    assign layer_0[6993] = in[585]; 
    assign layer_0[6994] = in[298] & in[693]; 
    assign layer_0[6995] = in[584]; 
    assign layer_0[6996] = in[444]; 
    assign layer_0[6997] = ~in[623] | (in[623] & in[617]); 
    assign layer_0[6998] = ~(in[286] ^ in[41]); 
    assign layer_0[6999] = ~(in[579] | in[693]); 
    assign layer_0[7000] = in[111] & in[13]; 
    assign layer_0[7001] = ~in[650]; 
    assign layer_0[7002] = in[519] | in[268]; 
    assign layer_0[7003] = ~(in[225] ^ in[731]); 
    assign layer_0[7004] = ~(in[584] ^ in[586]); 
    assign layer_0[7005] = ~in[161]; 
    assign layer_0[7006] = in[459] ^ in[311]; 
    assign layer_0[7007] = ~(in[342] | in[297]); 
    assign layer_0[7008] = in[458] & in[339]; 
    assign layer_0[7009] = in[728] ^ in[699]; 
    assign layer_0[7010] = in[247] ^ in[378]; 
    assign layer_0[7011] = ~(in[383] | in[96]); 
    assign layer_0[7012] = in[489] & ~in[466]; 
    assign layer_0[7013] = in[483] & ~in[379]; 
    assign layer_0[7014] = in[600] ^ in[487]; 
    assign layer_0[7015] = in[8]; 
    assign layer_0[7016] = in[419] | in[120]; 
    assign layer_0[7017] = in[254]; 
    assign layer_0[7018] = ~in[643] | (in[643] & in[740]); 
    assign layer_0[7019] = ~(in[474] ^ in[688]); 
    assign layer_0[7020] = in[222] ^ in[219]; 
    assign layer_0[7021] = ~(in[551] ^ in[86]); 
    assign layer_0[7022] = in[367] & ~in[659]; 
    assign layer_0[7023] = ~(in[487] ^ in[619]); 
    assign layer_0[7024] = in[675] & in[670]; 
    assign layer_0[7025] = ~in[280] | (in[280] & in[240]); 
    assign layer_0[7026] = in[66]; 
    assign layer_0[7027] = in[176]; 
    assign layer_0[7028] = in[745] | in[609]; 
    assign layer_0[7029] = in[361] & ~in[659]; 
    assign layer_0[7030] = in[99] & ~in[705]; 
    assign layer_0[7031] = in[626] & ~in[468]; 
    assign layer_0[7032] = ~in[90]; 
    assign layer_0[7033] = in[372] & ~in[759]; 
    assign layer_0[7034] = ~(in[372] ^ in[198]); 
    assign layer_0[7035] = ~in[198]; 
    assign layer_0[7036] = in[146] & ~in[737]; 
    assign layer_0[7037] = ~in[673] | (in[756] & in[673]); 
    assign layer_0[7038] = in[383] | in[467]; 
    assign layer_0[7039] = ~in[738]; 
    assign layer_0[7040] = ~(in[429] & in[94]); 
    assign layer_0[7041] = in[53] & ~in[31]; 
    assign layer_0[7042] = in[296] & ~in[346]; 
    assign layer_0[7043] = ~(in[661] | in[57]); 
    assign layer_0[7044] = in[598] ^ in[301]; 
    assign layer_0[7045] = ~(in[50] ^ in[299]); 
    assign layer_0[7046] = ~(in[142] | in[666]); 
    assign layer_0[7047] = ~(in[203] ^ in[651]); 
    assign layer_0[7048] = in[630] | in[7]; 
    assign layer_0[7049] = ~(in[399] ^ in[300]); 
    assign layer_0[7050] = in[632] ^ in[641]; 
    assign layer_0[7051] = in[641] & in[99]; 
    assign layer_0[7052] = in[6] & in[733]; 
    assign layer_0[7053] = ~in[475] | (in[475] & in[715]); 
    assign layer_0[7054] = in[85] & in[206]; 
    assign layer_0[7055] = in[267] ^ in[595]; 
    assign layer_0[7056] = in[675]; 
    assign layer_0[7057] = in[115] & ~in[581]; 
    assign layer_0[7058] = in[617] & ~in[81]; 
    assign layer_0[7059] = ~(in[468] | in[609]); 
    assign layer_0[7060] = in[218]; 
    assign layer_0[7061] = ~(in[473] ^ in[599]); 
    assign layer_0[7062] = ~(in[423] ^ in[346]); 
    assign layer_0[7063] = in[503] & ~in[394]; 
    assign layer_0[7064] = in[310] & in[327]; 
    assign layer_0[7065] = in[10] | in[728]; 
    assign layer_0[7066] = in[23] & in[412]; 
    assign layer_0[7067] = in[376] & ~in[505]; 
    assign layer_0[7068] = ~(in[9] & in[222]); 
    assign layer_0[7069] = in[622]; 
    assign layer_0[7070] = in[26]; 
    assign layer_0[7071] = in[474] ^ in[472]; 
    assign layer_0[7072] = in[616]; 
    assign layer_0[7073] = ~(in[522] ^ in[713]); 
    assign layer_0[7074] = in[139] ^ in[656]; 
    assign layer_0[7075] = in[29] ^ in[712]; 
    assign layer_0[7076] = in[376]; 
    assign layer_0[7077] = in[748] & ~in[649]; 
    assign layer_0[7078] = in[712] & in[564]; 
    assign layer_0[7079] = in[276] & ~in[342]; 
    assign layer_0[7080] = in[697] ^ in[695]; 
    assign layer_0[7081] = ~in[21]; 
    assign layer_0[7082] = ~in[49]; 
    assign layer_0[7083] = ~(in[276] ^ in[435]); 
    assign layer_0[7084] = in[226] ^ in[50]; 
    assign layer_0[7085] = in[491] ^ in[488]; 
    assign layer_0[7086] = ~in[310] | (in[310] & in[570]); 
    assign layer_0[7087] = ~(in[734] ^ in[620]); 
    assign layer_0[7088] = 1'b0; 
    assign layer_0[7089] = in[69]; 
    assign layer_0[7090] = ~(in[709] | in[541]); 
    assign layer_0[7091] = in[396] & ~in[692]; 
    assign layer_0[7092] = ~(in[712] ^ in[209]); 
    assign layer_0[7093] = in[108] ^ in[316]; 
    assign layer_0[7094] = ~(in[677] | in[224]); 
    assign layer_0[7095] = ~(in[430] ^ in[476]); 
    assign layer_0[7096] = ~in[598]; 
    assign layer_0[7097] = in[633]; 
    assign layer_0[7098] = in[341] & ~in[602]; 
    assign layer_0[7099] = in[659] & ~in[648]; 
    assign layer_0[7100] = in[560] | in[442]; 
    assign layer_0[7101] = ~in[757] | (in[757] & in[767]); 
    assign layer_0[7102] = in[423] & ~in[387]; 
    assign layer_0[7103] = ~(in[653] & in[338]); 
    assign layer_0[7104] = ~in[179] | (in[724] & in[179]); 
    assign layer_0[7105] = in[448] & in[660]; 
    assign layer_0[7106] = ~(in[299] ^ in[520]); 
    assign layer_0[7107] = in[411] & in[684]; 
    assign layer_0[7108] = ~(in[540] & in[482]); 
    assign layer_0[7109] = in[603] ^ in[178]; 
    assign layer_0[7110] = in[576] & ~in[429]; 
    assign layer_0[7111] = in[684] ^ in[206]; 
    assign layer_0[7112] = in[596] ^ in[662]; 
    assign layer_0[7113] = ~(in[135] & in[156]); 
    assign layer_0[7114] = ~(in[283] ^ in[142]); 
    assign layer_0[7115] = in[349] | in[287]; 
    assign layer_0[7116] = ~(in[364] ^ in[654]); 
    assign layer_0[7117] = in[645] ^ in[476]; 
    assign layer_0[7118] = ~in[566] | (in[566] & in[286]); 
    assign layer_0[7119] = in[461] & in[316]; 
    assign layer_0[7120] = ~(in[363] & in[603]); 
    assign layer_0[7121] = in[707] ^ in[717]; 
    assign layer_0[7122] = in[641] ^ in[97]; 
    assign layer_0[7123] = in[129] ^ in[130]; 
    assign layer_0[7124] = ~in[41]; 
    assign layer_0[7125] = ~(in[34] & in[254]); 
    assign layer_0[7126] = ~in[613] | (in[619] & in[613]); 
    assign layer_0[7127] = ~(in[529] | in[533]); 
    assign layer_0[7128] = ~in[263] | (in[263] & in[312]); 
    assign layer_0[7129] = in[520] & ~in[211]; 
    assign layer_0[7130] = in[534]; 
    assign layer_0[7131] = in[532] ^ in[60]; 
    assign layer_0[7132] = in[404] & ~in[731]; 
    assign layer_0[7133] = ~(in[490] & in[601]); 
    assign layer_0[7134] = in[356] ^ in[420]; 
    assign layer_0[7135] = ~(in[437] ^ in[80]); 
    assign layer_0[7136] = in[382] & ~in[605]; 
    assign layer_0[7137] = in[583] ^ in[662]; 
    assign layer_0[7138] = in[647] & in[549]; 
    assign layer_0[7139] = ~(in[760] ^ in[731]); 
    assign layer_0[7140] = ~(in[231] | in[314]); 
    assign layer_0[7141] = ~(in[352] ^ in[45]); 
    assign layer_0[7142] = in[286] & ~in[274]; 
    assign layer_0[7143] = ~(in[674] ^ in[34]); 
    assign layer_0[7144] = ~in[128]; 
    assign layer_0[7145] = ~in[487] | (in[487] & in[493]); 
    assign layer_0[7146] = ~(in[39] ^ in[556]); 
    assign layer_0[7147] = ~in[230]; 
    assign layer_0[7148] = in[160] ^ in[506]; 
    assign layer_0[7149] = in[617] | in[601]; 
    assign layer_0[7150] = ~(in[347] ^ in[218]); 
    assign layer_0[7151] = in[470] & in[90]; 
    assign layer_0[7152] = ~in[147] | (in[339] & in[147]); 
    assign layer_0[7153] = ~in[156] | (in[156] & in[616]); 
    assign layer_0[7154] = ~(in[581] | in[586]); 
    assign layer_0[7155] = ~in[551]; 
    assign layer_0[7156] = in[520] | in[46]; 
    assign layer_0[7157] = ~(in[104] & in[614]); 
    assign layer_0[7158] = in[725] & ~in[3]; 
    assign layer_0[7159] = ~(in[463] ^ in[79]); 
    assign layer_0[7160] = ~(in[699] ^ in[282]); 
    assign layer_0[7161] = ~(in[323] | in[623]); 
    assign layer_0[7162] = in[130] | in[766]; 
    assign layer_0[7163] = ~(in[221] | in[746]); 
    assign layer_0[7164] = ~in[248] | (in[248] & in[177]); 
    assign layer_0[7165] = ~in[302]; 
    assign layer_0[7166] = in[319] ^ in[300]; 
    assign layer_0[7167] = ~(in[657] ^ in[673]); 
    assign layer_0[7168] = in[536] ^ in[283]; 
    assign layer_0[7169] = in[615] ^ in[566]; 
    assign layer_0[7170] = in[172] & ~in[259]; 
    assign layer_0[7171] = ~(in[685] ^ in[471]); 
    assign layer_0[7172] = in[326] & ~in[278]; 
    assign layer_0[7173] = in[341] ^ in[143]; 
    assign layer_0[7174] = in[44] & ~in[30]; 
    assign layer_0[7175] = in[644] & ~in[740]; 
    assign layer_0[7176] = in[130] ^ in[550]; 
    assign layer_0[7177] = in[456] & ~in[275]; 
    assign layer_0[7178] = in[622] ^ in[625]; 
    assign layer_0[7179] = in[200] & ~in[714]; 
    assign layer_0[7180] = ~in[607] | (in[712] & in[607]); 
    assign layer_0[7181] = in[183] & ~in[320]; 
    assign layer_0[7182] = ~(in[640] ^ in[619]); 
    assign layer_0[7183] = in[99]; 
    assign layer_0[7184] = in[502] & ~in[493]; 
    assign layer_0[7185] = in[289] & ~in[636]; 
    assign layer_0[7186] = ~(in[673] ^ in[691]); 
    assign layer_0[7187] = ~in[277] | (in[681] & in[277]); 
    assign layer_0[7188] = in[140] & ~in[261]; 
    assign layer_0[7189] = in[228] ^ in[46]; 
    assign layer_0[7190] = in[125] | in[157]; 
    assign layer_0[7191] = ~in[286]; 
    assign layer_0[7192] = ~in[96] | (in[96] & in[547]); 
    assign layer_0[7193] = ~in[263] | (in[749] & in[263]); 
    assign layer_0[7194] = in[753] & ~in[619]; 
    assign layer_0[7195] = in[712]; 
    assign layer_0[7196] = ~(in[614] ^ in[235]); 
    assign layer_0[7197] = ~(in[19] & in[292]); 
    assign layer_0[7198] = ~in[536]; 
    assign layer_0[7199] = in[35] & ~in[587]; 
    assign layer_0[7200] = ~(in[644] ^ in[712]); 
    assign layer_0[7201] = ~(in[680] & in[278]); 
    assign layer_0[7202] = in[712] ^ in[692]; 
    assign layer_0[7203] = in[618]; 
    assign layer_0[7204] = ~(in[586] | in[299]); 
    assign layer_0[7205] = in[491] ^ in[157]; 
    assign layer_0[7206] = ~in[276] | (in[551] & in[276]); 
    assign layer_0[7207] = 1'b0; 
    assign layer_0[7208] = ~(in[648] ^ in[469]); 
    assign layer_0[7209] = in[45] ^ in[698]; 
    assign layer_0[7210] = ~in[580]; 
    assign layer_0[7211] = in[313] & ~in[643]; 
    assign layer_0[7212] = ~(in[756] & in[231]); 
    assign layer_0[7213] = in[336] ^ in[342]; 
    assign layer_0[7214] = in[586] & ~in[592]; 
    assign layer_0[7215] = in[296] ^ in[109]; 
    assign layer_0[7216] = ~in[327] | (in[327] & in[58]); 
    assign layer_0[7217] = in[750] | in[647]; 
    assign layer_0[7218] = ~(in[321] ^ in[392]); 
    assign layer_0[7219] = in[179] ^ in[520]; 
    assign layer_0[7220] = ~in[377]; 
    assign layer_0[7221] = in[228] | in[478]; 
    assign layer_0[7222] = ~in[589] | (in[589] & in[488]); 
    assign layer_0[7223] = in[507] | in[113]; 
    assign layer_0[7224] = ~(in[129] ^ in[157]); 
    assign layer_0[7225] = in[491] ^ in[345]; 
    assign layer_0[7226] = ~in[135] | (in[135] & in[643]); 
    assign layer_0[7227] = ~(in[542] ^ in[405]); 
    assign layer_0[7228] = ~(in[654] | in[605]); 
    assign layer_0[7229] = in[489] | in[63]; 
    assign layer_0[7230] = ~(in[66] ^ in[751]); 
    assign layer_0[7231] = ~(in[714] ^ in[618]); 
    assign layer_0[7232] = in[51]; 
    assign layer_0[7233] = ~(in[92] ^ in[356]); 
    assign layer_0[7234] = in[617] & ~in[355]; 
    assign layer_0[7235] = ~(in[348] ^ in[203]); 
    assign layer_0[7236] = in[584]; 
    assign layer_0[7237] = ~(in[242] | in[319]); 
    assign layer_0[7238] = ~in[390] | (in[390] & in[662]); 
    assign layer_0[7239] = in[474] & ~in[271]; 
    assign layer_0[7240] = ~in[727] | (in[727] & in[493]); 
    assign layer_0[7241] = in[78] ^ in[478]; 
    assign layer_0[7242] = ~in[692] | (in[173] & in[692]); 
    assign layer_0[7243] = ~(in[648] & in[692]); 
    assign layer_0[7244] = in[233] ^ in[52]; 
    assign layer_0[7245] = ~(in[581] | in[591]); 
    assign layer_0[7246] = in[732] & in[745]; 
    assign layer_0[7247] = ~in[91] | (in[243] & in[91]); 
    assign layer_0[7248] = in[99] & ~in[44]; 
    assign layer_0[7249] = ~(in[621] ^ in[129]); 
    assign layer_0[7250] = in[553] ^ in[611]; 
    assign layer_0[7251] = ~(in[372] ^ in[765]); 
    assign layer_0[7252] = in[392] & ~in[628]; 
    assign layer_0[7253] = ~(in[477] & in[327]); 
    assign layer_0[7254] = in[190] | in[540]; 
    assign layer_0[7255] = ~(in[92] & in[360]); 
    assign layer_0[7256] = in[586] & ~in[693]; 
    assign layer_0[7257] = ~(in[682] | in[244]); 
    assign layer_0[7258] = in[536] ^ in[600]; 
    assign layer_0[7259] = ~(in[572] ^ in[665]); 
    assign layer_0[7260] = in[152] & ~in[349]; 
    assign layer_0[7261] = ~in[463]; 
    assign layer_0[7262] = ~(in[361] ^ in[706]); 
    assign layer_0[7263] = in[172]; 
    assign layer_0[7264] = in[459] & in[344]; 
    assign layer_0[7265] = in[600]; 
    assign layer_0[7266] = ~in[659]; 
    assign layer_0[7267] = ~(in[657] ^ in[675]); 
    assign layer_0[7268] = in[684] ^ in[614]; 
    assign layer_0[7269] = ~(in[273] & in[639]); 
    assign layer_0[7270] = in[520] ^ in[521]; 
    assign layer_0[7271] = ~in[24]; 
    assign layer_0[7272] = in[24]; 
    assign layer_0[7273] = in[550] | in[500]; 
    assign layer_0[7274] = ~(in[294] | in[7]); 
    assign layer_0[7275] = in[206] & in[377]; 
    assign layer_0[7276] = in[65]; 
    assign layer_0[7277] = in[372] & ~in[340]; 
    assign layer_0[7278] = in[655] | in[759]; 
    assign layer_0[7279] = in[372] ^ in[747]; 
    assign layer_0[7280] = in[743]; 
    assign layer_0[7281] = in[365] & ~in[697]; 
    assign layer_0[7282] = ~(in[108] | in[50]); 
    assign layer_0[7283] = ~(in[363] ^ in[475]); 
    assign layer_0[7284] = ~(in[442] & in[282]); 
    assign layer_0[7285] = ~(in[417] & in[62]); 
    assign layer_0[7286] = ~(in[372] ^ in[265]); 
    assign layer_0[7287] = ~in[588]; 
    assign layer_0[7288] = ~(in[475] | in[668]); 
    assign layer_0[7289] = ~in[547]; 
    assign layer_0[7290] = in[603] & ~in[160]; 
    assign layer_0[7291] = ~in[18] | (in[18] & in[452]); 
    assign layer_0[7292] = in[72] ^ in[356]; 
    assign layer_0[7293] = in[347] ^ in[62]; 
    assign layer_0[7294] = in[408] & in[548]; 
    assign layer_0[7295] = ~in[710]; 
    assign layer_0[7296] = ~in[650] | (in[650] & in[494]); 
    assign layer_0[7297] = ~(in[263] | in[16]); 
    assign layer_0[7298] = in[664]; 
    assign layer_0[7299] = ~(in[413] ^ in[102]); 
    assign layer_0[7300] = ~in[661]; 
    assign layer_0[7301] = in[696] ^ in[747]; 
    assign layer_0[7302] = in[634] ^ in[76]; 
    assign layer_0[7303] = in[695] ^ in[279]; 
    assign layer_0[7304] = ~in[582]; 
    assign layer_0[7305] = ~in[506]; 
    assign layer_0[7306] = in[654]; 
    assign layer_0[7307] = ~(in[611] ^ in[652]); 
    assign layer_0[7308] = ~in[144]; 
    assign layer_0[7309] = in[468] ^ in[462]; 
    assign layer_0[7310] = ~(in[519] | in[467]); 
    assign layer_0[7311] = in[487] & ~in[324]; 
    assign layer_0[7312] = ~in[468] | (in[468] & in[311]); 
    assign layer_0[7313] = in[158] ^ in[49]; 
    assign layer_0[7314] = ~in[107] | (in[107] & in[520]); 
    assign layer_0[7315] = in[412] | in[66]; 
    assign layer_0[7316] = ~(in[483] ^ in[748]); 
    assign layer_0[7317] = ~(in[0] | in[696]); 
    assign layer_0[7318] = in[605] & in[527]; 
    assign layer_0[7319] = ~in[678]; 
    assign layer_0[7320] = ~in[20] | (in[20] & in[652]); 
    assign layer_0[7321] = in[265] & ~in[536]; 
    assign layer_0[7322] = ~(in[614] ^ in[600]); 
    assign layer_0[7323] = in[467] ^ in[297]; 
    assign layer_0[7324] = in[298] ^ in[386]; 
    assign layer_0[7325] = in[267] & ~in[681]; 
    assign layer_0[7326] = in[382]; 
    assign layer_0[7327] = in[132] & ~in[758]; 
    assign layer_0[7328] = in[442] ^ in[178]; 
    assign layer_0[7329] = ~(in[393] & in[182]); 
    assign layer_0[7330] = in[691] ^ in[676]; 
    assign layer_0[7331] = in[694] & ~in[621]; 
    assign layer_0[7332] = in[660] & in[113]; 
    assign layer_0[7333] = ~in[266] | (in[266] & in[728]); 
    assign layer_0[7334] = in[324]; 
    assign layer_0[7335] = ~(in[56] & in[759]); 
    assign layer_0[7336] = in[83] & in[340]; 
    assign layer_0[7337] = ~(in[340] | in[34]); 
    assign layer_0[7338] = in[387] | in[322]; 
    assign layer_0[7339] = in[757] ^ in[658]; 
    assign layer_0[7340] = ~(in[112] & in[589]); 
    assign layer_0[7341] = ~in[248]; 
    assign layer_0[7342] = ~in[92]; 
    assign layer_0[7343] = in[22]; 
    assign layer_0[7344] = ~(in[706] | in[267]); 
    assign layer_0[7345] = in[129] & ~in[312]; 
    assign layer_0[7346] = ~(in[67] | in[698]); 
    assign layer_0[7347] = in[49] ^ in[474]; 
    assign layer_0[7348] = ~(in[391] & in[394]); 
    assign layer_0[7349] = 1'b1; 
    assign layer_0[7350] = ~(in[324] ^ in[618]); 
    assign layer_0[7351] = in[680] & ~in[589]; 
    assign layer_0[7352] = in[634] & ~in[725]; 
    assign layer_0[7353] = ~in[491] | (in[516] & in[491]); 
    assign layer_0[7354] = ~in[6] | (in[6] & in[261]); 
    assign layer_0[7355] = ~in[519] | (in[519] & in[652]); 
    assign layer_0[7356] = in[401] & in[111]; 
    assign layer_0[7357] = ~in[709] | (in[582] & in[709]); 
    assign layer_0[7358] = in[49]; 
    assign layer_0[7359] = in[697] | in[666]; 
    assign layer_0[7360] = in[73] ^ in[93]; 
    assign layer_0[7361] = in[554] ^ in[555]; 
    assign layer_0[7362] = in[235] & ~in[19]; 
    assign layer_0[7363] = in[138]; 
    assign layer_0[7364] = ~in[572]; 
    assign layer_0[7365] = in[412] & ~in[613]; 
    assign layer_0[7366] = in[377] ^ in[211]; 
    assign layer_0[7367] = in[309] ^ in[340]; 
    assign layer_0[7368] = in[380] ^ in[253]; 
    assign layer_0[7369] = in[19]; 
    assign layer_0[7370] = in[435] | in[565]; 
    assign layer_0[7371] = ~in[713]; 
    assign layer_0[7372] = ~in[233] | (in[520] & in[233]); 
    assign layer_0[7373] = ~(in[95] ^ in[723]); 
    assign layer_0[7374] = in[711] & ~in[161]; 
    assign layer_0[7375] = in[570]; 
    assign layer_0[7376] = ~in[230]; 
    assign layer_0[7377] = ~(in[44] & in[519]); 
    assign layer_0[7378] = in[660] ^ in[397]; 
    assign layer_0[7379] = in[701] ^ in[635]; 
    assign layer_0[7380] = ~in[361] | (in[759] & in[361]); 
    assign layer_0[7381] = ~in[231] | (in[468] & in[231]); 
    assign layer_0[7382] = ~(in[399] ^ in[285]); 
    assign layer_0[7383] = ~(in[157] ^ in[371]); 
    assign layer_0[7384] = in[633]; 
    assign layer_0[7385] = ~(in[338] | in[239]); 
    assign layer_0[7386] = in[618] ^ in[554]; 
    assign layer_0[7387] = in[533] & ~in[483]; 
    assign layer_0[7388] = ~(in[735] | in[586]); 
    assign layer_0[7389] = in[562] ^ in[344]; 
    assign layer_0[7390] = in[332]; 
    assign layer_0[7391] = ~in[645]; 
    assign layer_0[7392] = ~in[483]; 
    assign layer_0[7393] = in[458] & ~in[305]; 
    assign layer_0[7394] = ~(in[645] ^ in[656]); 
    assign layer_0[7395] = ~(in[618] | in[585]); 
    assign layer_0[7396] = ~(in[589] ^ in[467]); 
    assign layer_0[7397] = ~in[108]; 
    assign layer_0[7398] = in[279] | in[725]; 
    assign layer_0[7399] = in[459]; 
    assign layer_0[7400] = in[114] & ~in[635]; 
    assign layer_0[7401] = in[231] & ~in[717]; 
    assign layer_0[7402] = ~in[580] | (in[748] & in[580]); 
    assign layer_0[7403] = ~(in[738] ^ in[744]); 
    assign layer_0[7404] = in[474] & in[757]; 
    assign layer_0[7405] = ~in[396] | (in[699] & in[396]); 
    assign layer_0[7406] = ~(in[149] & in[219]); 
    assign layer_0[7407] = in[121] | in[661]; 
    assign layer_0[7408] = in[196] ^ in[423]; 
    assign layer_0[7409] = ~in[61]; 
    assign layer_0[7410] = 1'b0; 
    assign layer_0[7411] = ~(in[604] | in[518]); 
    assign layer_0[7412] = ~in[403]; 
    assign layer_0[7413] = ~in[27]; 
    assign layer_0[7414] = in[301]; 
    assign layer_0[7415] = in[579] ^ in[723]; 
    assign layer_0[7416] = in[268] & ~in[162]; 
    assign layer_0[7417] = in[50] | in[675]; 
    assign layer_0[7418] = ~in[664] | (in[664] & in[543]); 
    assign layer_0[7419] = in[761] | in[697]; 
    assign layer_0[7420] = ~in[726] | (in[665] & in[726]); 
    assign layer_0[7421] = in[630] ^ in[283]; 
    assign layer_0[7422] = in[681]; 
    assign layer_0[7423] = ~(in[588] ^ in[590]); 
    assign layer_0[7424] = in[339] | in[692]; 
    assign layer_0[7425] = ~(in[331] & in[208]); 
    assign layer_0[7426] = ~in[528] | (in[273] & in[528]); 
    assign layer_0[7427] = in[111] & in[403]; 
    assign layer_0[7428] = ~(in[189] | in[537]); 
    assign layer_0[7429] = in[611] & ~in[606]; 
    assign layer_0[7430] = in[496]; 
    assign layer_0[7431] = ~in[745] | (in[629] & in[745]); 
    assign layer_0[7432] = in[760] | in[96]; 
    assign layer_0[7433] = ~in[504]; 
    assign layer_0[7434] = in[677] ^ in[585]; 
    assign layer_0[7435] = in[219] & ~in[762]; 
    assign layer_0[7436] = ~(in[74] ^ in[68]); 
    assign layer_0[7437] = ~(in[141] ^ in[237]); 
    assign layer_0[7438] = in[672] & ~in[42]; 
    assign layer_0[7439] = in[673]; 
    assign layer_0[7440] = in[678] | in[745]; 
    assign layer_0[7441] = ~(in[331] ^ in[693]); 
    assign layer_0[7442] = in[277] ^ in[722]; 
    assign layer_0[7443] = ~in[419] | (in[419] & in[99]); 
    assign layer_0[7444] = ~in[211] | (in[46] & in[211]); 
    assign layer_0[7445] = in[226] & in[8]; 
    assign layer_0[7446] = ~(in[79] & in[618]); 
    assign layer_0[7447] = ~(in[364] ^ in[94]); 
    assign layer_0[7448] = ~(in[631] | in[605]); 
    assign layer_0[7449] = in[263] | in[708]; 
    assign layer_0[7450] = ~(in[556] ^ in[266]); 
    assign layer_0[7451] = in[204] & ~in[557]; 
    assign layer_0[7452] = in[299]; 
    assign layer_0[7453] = in[89] & in[615]; 
    assign layer_0[7454] = in[746] ^ in[698]; 
    assign layer_0[7455] = ~(in[670] & in[665]); 
    assign layer_0[7456] = ~(in[45] ^ in[681]); 
    assign layer_0[7457] = in[742] ^ in[744]; 
    assign layer_0[7458] = in[710] & ~in[83]; 
    assign layer_0[7459] = ~in[329]; 
    assign layer_0[7460] = in[29] ^ in[752]; 
    assign layer_0[7461] = in[615] ^ in[630]; 
    assign layer_0[7462] = in[759] & ~in[681]; 
    assign layer_0[7463] = in[137] ^ in[680]; 
    assign layer_0[7464] = ~in[124]; 
    assign layer_0[7465] = in[312] ^ in[68]; 
    assign layer_0[7466] = ~(in[571] ^ in[666]); 
    assign layer_0[7467] = ~(in[127] | in[705]); 
    assign layer_0[7468] = in[642] ^ in[28]; 
    assign layer_0[7469] = in[299] ^ in[346]; 
    assign layer_0[7470] = in[278] | in[524]; 
    assign layer_0[7471] = ~in[217]; 
    assign layer_0[7472] = in[318] ^ in[670]; 
    assign layer_0[7473] = in[671]; 
    assign layer_0[7474] = ~(in[378] ^ in[411]); 
    assign layer_0[7475] = ~(in[440] & in[408]); 
    assign layer_0[7476] = in[371] ^ in[396]; 
    assign layer_0[7477] = ~(in[220] ^ in[236]); 
    assign layer_0[7478] = ~(in[680] ^ in[211]); 
    assign layer_0[7479] = ~(in[389] | in[168]); 
    assign layer_0[7480] = in[145] ^ in[350]; 
    assign layer_0[7481] = in[618]; 
    assign layer_0[7482] = in[427] & ~in[715]; 
    assign layer_0[7483] = ~(in[30] ^ in[347]); 
    assign layer_0[7484] = in[190]; 
    assign layer_0[7485] = ~(in[594] ^ in[445]); 
    assign layer_0[7486] = ~in[509]; 
    assign layer_0[7487] = in[595] & ~in[396]; 
    assign layer_0[7488] = in[595] | in[28]; 
    assign layer_0[7489] = in[445]; 
    assign layer_0[7490] = ~in[710] | (in[146] & in[710]); 
    assign layer_0[7491] = ~in[308] | (in[308] & in[342]); 
    assign layer_0[7492] = in[338]; 
    assign layer_0[7493] = ~(in[458] & in[457]); 
    assign layer_0[7494] = in[363] ^ in[470]; 
    assign layer_0[7495] = in[657] & in[599]; 
    assign layer_0[7496] = in[21] | in[527]; 
    assign layer_0[7497] = in[724] ^ in[25]; 
    assign layer_0[7498] = in[738] & ~in[631]; 
    assign layer_0[7499] = ~in[487] | (in[487] & in[265]); 
    assign layer_0[7500] = in[29] & ~in[635]; 
    assign layer_0[7501] = ~(in[638] ^ in[85]); 
    assign layer_0[7502] = in[420] & ~in[92]; 
    assign layer_0[7503] = ~(in[412] & in[230]); 
    assign layer_0[7504] = in[600] ^ in[604]; 
    assign layer_0[7505] = in[54] ^ in[208]; 
    assign layer_0[7506] = in[140] & in[8]; 
    assign layer_0[7507] = ~in[560] | (in[560] & in[683]); 
    assign layer_0[7508] = ~in[243] | (in[665] & in[243]); 
    assign layer_0[7509] = ~(in[522] & in[474]); 
    assign layer_0[7510] = ~(in[552] ^ in[13]); 
    assign layer_0[7511] = ~(in[554] ^ in[758]); 
    assign layer_0[7512] = in[691] ^ in[747]; 
    assign layer_0[7513] = ~in[719] | (in[719] & in[402]); 
    assign layer_0[7514] = ~in[411]; 
    assign layer_0[7515] = in[296] | in[297]; 
    assign layer_0[7516] = ~(in[664] | in[647]); 
    assign layer_0[7517] = ~(in[339] & in[680]); 
    assign layer_0[7518] = ~(in[498] ^ in[616]); 
    assign layer_0[7519] = in[157] ^ in[680]; 
    assign layer_0[7520] = in[479] & in[391]; 
    assign layer_0[7521] = ~(in[637] | in[307]); 
    assign layer_0[7522] = ~(in[615] ^ in[471]); 
    assign layer_0[7523] = ~(in[183] | in[340]); 
    assign layer_0[7524] = in[615] & in[10]; 
    assign layer_0[7525] = ~(in[265] | in[381]); 
    assign layer_0[7526] = ~(in[596] | in[763]); 
    assign layer_0[7527] = in[34] ^ in[555]; 
    assign layer_0[7528] = in[430] & ~in[48]; 
    assign layer_0[7529] = ~(in[430] ^ in[587]); 
    assign layer_0[7530] = in[354]; 
    assign layer_0[7531] = ~(in[380] ^ in[264]); 
    assign layer_0[7532] = ~(in[91] ^ in[281]); 
    assign layer_0[7533] = in[292] | in[724]; 
    assign layer_0[7534] = in[248] ^ in[692]; 
    assign layer_0[7535] = in[13] ^ in[95]; 
    assign layer_0[7536] = ~(in[586] | in[99]); 
    assign layer_0[7537] = ~(in[399] | in[723]); 
    assign layer_0[7538] = ~(in[745] ^ in[714]); 
    assign layer_0[7539] = in[473] ^ in[470]; 
    assign layer_0[7540] = in[406] & in[310]; 
    assign layer_0[7541] = in[691] & ~in[267]; 
    assign layer_0[7542] = in[435]; 
    assign layer_0[7543] = in[327]; 
    assign layer_0[7544] = 1'b0; 
    assign layer_0[7545] = ~(in[239] ^ in[110]); 
    assign layer_0[7546] = ~in[584] | (in[584] & in[504]); 
    assign layer_0[7547] = in[110]; 
    assign layer_0[7548] = in[693] & ~in[600]; 
    assign layer_0[7549] = ~in[298] | (in[370] & in[298]); 
    assign layer_0[7550] = ~in[480] | (in[480] & in[493]); 
    assign layer_0[7551] = ~(in[295] & in[66]); 
    assign layer_0[7552] = ~(in[565] ^ in[297]); 
    assign layer_0[7553] = in[655]; 
    assign layer_0[7554] = ~in[415] | (in[415] & in[734]); 
    assign layer_0[7555] = ~(in[731] ^ in[586]); 
    assign layer_0[7556] = in[556] | in[208]; 
    assign layer_0[7557] = ~(in[323] ^ in[271]); 
    assign layer_0[7558] = in[388] ^ in[14]; 
    assign layer_0[7559] = in[232] | in[38]; 
    assign layer_0[7560] = ~in[77] | (in[551] & in[77]); 
    assign layer_0[7561] = in[602] & ~in[730]; 
    assign layer_0[7562] = ~in[83]; 
    assign layer_0[7563] = in[654] & ~in[612]; 
    assign layer_0[7564] = ~(in[424] ^ in[345]); 
    assign layer_0[7565] = ~(in[750] | in[394]); 
    assign layer_0[7566] = in[227]; 
    assign layer_0[7567] = in[542] ^ in[272]; 
    assign layer_0[7568] = ~(in[572] ^ in[749]); 
    assign layer_0[7569] = in[462]; 
    assign layer_0[7570] = in[461] & ~in[95]; 
    assign layer_0[7571] = in[521] ^ in[254]; 
    assign layer_0[7572] = ~(in[163] ^ in[468]); 
    assign layer_0[7573] = ~in[475] | (in[688] & in[475]); 
    assign layer_0[7574] = ~(in[752] ^ in[223]); 
    assign layer_0[7575] = ~in[425]; 
    assign layer_0[7576] = ~in[746] | (in[746] & in[177]); 
    assign layer_0[7577] = in[632] ^ in[227]; 
    assign layer_0[7578] = ~in[242] | (in[45] & in[242]); 
    assign layer_0[7579] = ~(in[742] ^ in[661]); 
    assign layer_0[7580] = in[422] & ~in[539]; 
    assign layer_0[7581] = ~(in[70] & in[19]); 
    assign layer_0[7582] = in[45] & ~in[237]; 
    assign layer_0[7583] = ~in[279]; 
    assign layer_0[7584] = in[52]; 
    assign layer_0[7585] = ~(in[8] | in[447]); 
    assign layer_0[7586] = ~(in[462] | in[443]); 
    assign layer_0[7587] = in[265] & in[262]; 
    assign layer_0[7588] = in[626] ^ in[63]; 
    assign layer_0[7589] = in[84] | in[599]; 
    assign layer_0[7590] = in[387] ^ in[547]; 
    assign layer_0[7591] = ~(in[355] & in[110]); 
    assign layer_0[7592] = ~in[637] | (in[504] & in[637]); 
    assign layer_0[7593] = in[564] | in[682]; 
    assign layer_0[7594] = in[597] ^ in[602]; 
    assign layer_0[7595] = ~in[327]; 
    assign layer_0[7596] = ~(in[367] & in[153]); 
    assign layer_0[7597] = in[691] | in[355]; 
    assign layer_0[7598] = in[120]; 
    assign layer_0[7599] = ~(in[232] & in[713]); 
    assign layer_0[7600] = 1'b1; 
    assign layer_0[7601] = ~(in[255] | in[362]); 
    assign layer_0[7602] = in[407] & ~in[641]; 
    assign layer_0[7603] = in[565] ^ in[629]; 
    assign layer_0[7604] = ~in[380] | (in[62] & in[380]); 
    assign layer_0[7605] = in[326] & ~in[603]; 
    assign layer_0[7606] = in[618] ^ in[586]; 
    assign layer_0[7607] = in[622]; 
    assign layer_0[7608] = in[348] & ~in[597]; 
    assign layer_0[7609] = ~in[314]; 
    assign layer_0[7610] = ~(in[609] ^ in[505]); 
    assign layer_0[7611] = ~in[266]; 
    assign layer_0[7612] = 1'b0; 
    assign layer_0[7613] = ~in[591] | (in[591] & in[637]); 
    assign layer_0[7614] = in[614] & ~in[547]; 
    assign layer_0[7615] = in[629] ^ in[696]; 
    assign layer_0[7616] = ~in[211]; 
    assign layer_0[7617] = ~(in[553] ^ in[677]); 
    assign layer_0[7618] = in[242] & ~in[193]; 
    assign layer_0[7619] = in[725] | in[617]; 
    assign layer_0[7620] = in[279]; 
    assign layer_0[7621] = in[604]; 
    assign layer_0[7622] = ~in[355] | (in[242] & in[355]); 
    assign layer_0[7623] = ~in[218] | (in[218] & in[534]); 
    assign layer_0[7624] = ~(in[664] ^ in[712]); 
    assign layer_0[7625] = in[554] | in[698]; 
    assign layer_0[7626] = in[633] & ~in[708]; 
    assign layer_0[7627] = ~in[203] | (in[203] & in[47]); 
    assign layer_0[7628] = ~(in[221] | in[568]); 
    assign layer_0[7629] = in[740] ^ in[396]; 
    assign layer_0[7630] = ~(in[34] | in[733]); 
    assign layer_0[7631] = ~(in[68] ^ in[670]); 
    assign layer_0[7632] = in[231]; 
    assign layer_0[7633] = in[252] & ~in[738]; 
    assign layer_0[7634] = ~(in[460] | in[95]); 
    assign layer_0[7635] = in[631] ^ in[700]; 
    assign layer_0[7636] = in[458] ^ in[744]; 
    assign layer_0[7637] = in[192] | in[433]; 
    assign layer_0[7638] = in[397] ^ in[331]; 
    assign layer_0[7639] = ~(in[78] ^ in[395]); 
    assign layer_0[7640] = ~in[309]; 
    assign layer_0[7641] = ~in[202] | (in[202] & in[600]); 
    assign layer_0[7642] = in[750] ^ in[110]; 
    assign layer_0[7643] = ~in[195]; 
    assign layer_0[7644] = ~(in[646] ^ in[177]); 
    assign layer_0[7645] = ~(in[297] ^ in[652]); 
    assign layer_0[7646] = in[538] & in[378]; 
    assign layer_0[7647] = ~(in[308] & in[695]); 
    assign layer_0[7648] = ~in[699]; 
    assign layer_0[7649] = ~(in[552] ^ in[760]); 
    assign layer_0[7650] = ~(in[343] ^ in[66]); 
    assign layer_0[7651] = in[417] ^ in[38]; 
    assign layer_0[7652] = in[82] & in[365]; 
    assign layer_0[7653] = ~in[428]; 
    assign layer_0[7654] = ~in[317]; 
    assign layer_0[7655] = 1'b0; 
    assign layer_0[7656] = ~(in[432] ^ in[694]); 
    assign layer_0[7657] = ~(in[477] ^ in[242]); 
    assign layer_0[7658] = in[263] & ~in[563]; 
    assign layer_0[7659] = ~(in[462] | in[570]); 
    assign layer_0[7660] = ~in[94]; 
    assign layer_0[7661] = in[662] ^ in[476]; 
    assign layer_0[7662] = in[140] & ~in[552]; 
    assign layer_0[7663] = in[312] ^ in[520]; 
    assign layer_0[7664] = in[221] & ~in[246]; 
    assign layer_0[7665] = in[78] & ~in[247]; 
    assign layer_0[7666] = in[203] ^ in[357]; 
    assign layer_0[7667] = 1'b0; 
    assign layer_0[7668] = 1'b0; 
    assign layer_0[7669] = in[680] & ~in[600]; 
    assign layer_0[7670] = ~(in[516] & in[347]); 
    assign layer_0[7671] = in[664] & ~in[502]; 
    assign layer_0[7672] = ~in[19] | (in[679] & in[19]); 
    assign layer_0[7673] = ~in[325] | (in[586] & in[325]); 
    assign layer_0[7674] = ~in[724]; 
    assign layer_0[7675] = ~in[408] | (in[237] & in[408]); 
    assign layer_0[7676] = in[422] & in[660]; 
    assign layer_0[7677] = in[660] | in[719]; 
    assign layer_0[7678] = in[254] & in[82]; 
    assign layer_0[7679] = ~(in[634] & in[681]); 
    assign layer_0[7680] = in[474] & ~in[595]; 
    assign layer_0[7681] = in[162] & in[630]; 
    assign layer_0[7682] = in[448] ^ in[91]; 
    assign layer_0[7683] = ~(in[176] ^ in[249]); 
    assign layer_0[7684] = in[651] ^ in[579]; 
    assign layer_0[7685] = ~in[587]; 
    assign layer_0[7686] = in[534] | in[276]; 
    assign layer_0[7687] = ~(in[651] ^ in[587]); 
    assign layer_0[7688] = in[4] ^ in[635]; 
    assign layer_0[7689] = ~in[32] | (in[363] & in[32]); 
    assign layer_0[7690] = ~in[620] | (in[620] & in[457]); 
    assign layer_0[7691] = ~in[283] | (in[114] & in[283]); 
    assign layer_0[7692] = in[707]; 
    assign layer_0[7693] = ~(in[347] ^ in[330]); 
    assign layer_0[7694] = in[548] ^ in[205]; 
    assign layer_0[7695] = in[699] ^ in[315]; 
    assign layer_0[7696] = in[81] | in[466]; 
    assign layer_0[7697] = in[128] | in[327]; 
    assign layer_0[7698] = ~(in[520] ^ in[711]); 
    assign layer_0[7699] = in[402] ^ in[194]; 
    assign layer_0[7700] = ~(in[480] ^ in[305]); 
    assign layer_0[7701] = ~in[716] | (in[716] & in[745]); 
    assign layer_0[7702] = in[426] ^ in[404]; 
    assign layer_0[7703] = ~(in[252] ^ in[634]); 
    assign layer_0[7704] = ~(in[324] ^ in[345]); 
    assign layer_0[7705] = ~in[347] | (in[428] & in[347]); 
    assign layer_0[7706] = in[331] & ~in[619]; 
    assign layer_0[7707] = ~in[110] | (in[42] & in[110]); 
    assign layer_0[7708] = ~(in[30] ^ in[253]); 
    assign layer_0[7709] = in[706] ^ in[560]; 
    assign layer_0[7710] = ~in[457] | (in[650] & in[457]); 
    assign layer_0[7711] = ~in[666] | (in[225] & in[666]); 
    assign layer_0[7712] = ~(in[332] ^ in[454]); 
    assign layer_0[7713] = in[436] & in[45]; 
    assign layer_0[7714] = ~(in[614] & in[619]); 
    assign layer_0[7715] = in[460]; 
    assign layer_0[7716] = in[294] ^ in[46]; 
    assign layer_0[7717] = in[330] & in[602]; 
    assign layer_0[7718] = in[236] & in[488]; 
    assign layer_0[7719] = ~(in[364] ^ in[358]); 
    assign layer_0[7720] = ~(in[728] & in[746]); 
    assign layer_0[7721] = in[308]; 
    assign layer_0[7722] = ~in[160] | (in[160] & in[406]); 
    assign layer_0[7723] = in[672] ^ in[623]; 
    assign layer_0[7724] = in[681] & ~in[504]; 
    assign layer_0[7725] = ~(in[20] & in[234]); 
    assign layer_0[7726] = ~in[152] | (in[628] & in[152]); 
    assign layer_0[7727] = in[569] ^ in[652]; 
    assign layer_0[7728] = ~(in[141] | in[334]); 
    assign layer_0[7729] = ~in[265]; 
    assign layer_0[7730] = in[298]; 
    assign layer_0[7731] = in[727] ^ in[110]; 
    assign layer_0[7732] = ~(in[425] & in[312]); 
    assign layer_0[7733] = in[660] & ~in[296]; 
    assign layer_0[7734] = ~(in[716] | in[535]); 
    assign layer_0[7735] = in[440] & ~in[623]; 
    assign layer_0[7736] = ~in[277] | (in[277] & in[263]); 
    assign layer_0[7737] = in[327]; 
    assign layer_0[7738] = 1'b1; 
    assign layer_0[7739] = ~(in[580] ^ in[386]); 
    assign layer_0[7740] = ~in[93]; 
    assign layer_0[7741] = in[27] & ~in[225]; 
    assign layer_0[7742] = ~(in[531] | in[366]); 
    assign layer_0[7743] = ~in[712]; 
    assign layer_0[7744] = in[474] ^ in[19]; 
    assign layer_0[7745] = in[492] & in[283]; 
    assign layer_0[7746] = in[443] ^ in[741]; 
    assign layer_0[7747] = in[535]; 
    assign layer_0[7748] = in[712] & ~in[207]; 
    assign layer_0[7749] = in[110] | in[110]; 
    assign layer_0[7750] = ~(in[692] | in[716]); 
    assign layer_0[7751] = ~(in[660] ^ in[467]); 
    assign layer_0[7752] = in[118] ^ in[14]; 
    assign layer_0[7753] = in[36] & ~in[323]; 
    assign layer_0[7754] = in[694] ^ in[351]; 
    assign layer_0[7755] = ~in[728]; 
    assign layer_0[7756] = in[35] | in[113]; 
    assign layer_0[7757] = in[208] ^ in[179]; 
    assign layer_0[7758] = ~(in[586] ^ in[708]); 
    assign layer_0[7759] = ~in[646] | (in[646] & in[694]); 
    assign layer_0[7760] = 1'b1; 
    assign layer_0[7761] = ~in[644] | (in[644] & in[505]); 
    assign layer_0[7762] = ~(in[112] ^ in[211]); 
    assign layer_0[7763] = in[46] ^ in[111]; 
    assign layer_0[7764] = in[35]; 
    assign layer_0[7765] = ~in[466]; 
    assign layer_0[7766] = ~(in[56] & in[76]); 
    assign layer_0[7767] = ~(in[685] ^ in[308]); 
    assign layer_0[7768] = ~(in[226] ^ in[29]); 
    assign layer_0[7769] = in[411]; 
    assign layer_0[7770] = in[264] & ~in[55]; 
    assign layer_0[7771] = ~in[98]; 
    assign layer_0[7772] = in[613] | in[661]; 
    assign layer_0[7773] = ~(in[409] ^ in[570]); 
    assign layer_0[7774] = in[50] & in[316]; 
    assign layer_0[7775] = in[658]; 
    assign layer_0[7776] = in[239] ^ in[314]; 
    assign layer_0[7777] = ~(in[619] | in[411]); 
    assign layer_0[7778] = ~in[286] | (in[65] & in[286]); 
    assign layer_0[7779] = ~in[645] | (in[519] & in[645]); 
    assign layer_0[7780] = ~(in[418] | in[734]); 
    assign layer_0[7781] = ~(in[544] | in[82]); 
    assign layer_0[7782] = 1'b0; 
    assign layer_0[7783] = in[723] ^ in[597]; 
    assign layer_0[7784] = in[665] | in[628]; 
    assign layer_0[7785] = in[620] ^ in[40]; 
    assign layer_0[7786] = in[436]; 
    assign layer_0[7787] = in[645] | in[333]; 
    assign layer_0[7788] = in[725]; 
    assign layer_0[7789] = in[432] & in[517]; 
    assign layer_0[7790] = in[91] | in[491]; 
    assign layer_0[7791] = in[230] ^ in[700]; 
    assign layer_0[7792] = ~(in[128] ^ in[717]); 
    assign layer_0[7793] = ~(in[21] | in[615]); 
    assign layer_0[7794] = in[19] & in[323]; 
    assign layer_0[7795] = in[447] & ~in[54]; 
    assign layer_0[7796] = ~in[678] | (in[275] & in[678]); 
    assign layer_0[7797] = in[279] & ~in[182]; 
    assign layer_0[7798] = ~(in[221] & in[143]); 
    assign layer_0[7799] = in[733] | in[651]; 
    assign layer_0[7800] = in[241] & in[477]; 
    assign layer_0[7801] = ~in[714] | (in[128] & in[714]); 
    assign layer_0[7802] = ~(in[176] | in[242]); 
    assign layer_0[7803] = in[473] & ~in[557]; 
    assign layer_0[7804] = ~(in[298] ^ in[586]); 
    assign layer_0[7805] = in[424] ^ in[594]; 
    assign layer_0[7806] = ~(in[628] ^ in[615]); 
    assign layer_0[7807] = in[667] & ~in[125]; 
    assign layer_0[7808] = in[356] ^ in[342]; 
    assign layer_0[7809] = ~(in[450] & in[458]); 
    assign layer_0[7810] = in[150]; 
    assign layer_0[7811] = ~(in[744] ^ in[535]); 
    assign layer_0[7812] = in[281] & ~in[18]; 
    assign layer_0[7813] = ~in[554] | (in[554] & in[192]); 
    assign layer_0[7814] = ~in[425] | (in[425] & in[688]); 
    assign layer_0[7815] = in[599] & ~in[636]; 
    assign layer_0[7816] = ~(in[359] ^ in[322]); 
    assign layer_0[7817] = ~(in[662] ^ in[745]); 
    assign layer_0[7818] = in[56] & ~in[597]; 
    assign layer_0[7819] = in[446]; 
    assign layer_0[7820] = in[585] & in[616]; 
    assign layer_0[7821] = in[340] & ~in[726]; 
    assign layer_0[7822] = ~(in[243] & in[626]); 
    assign layer_0[7823] = in[266] ^ in[666]; 
    assign layer_0[7824] = ~(in[537] | in[534]); 
    assign layer_0[7825] = ~in[712]; 
    assign layer_0[7826] = ~(in[708] ^ in[494]); 
    assign layer_0[7827] = ~(in[93] | in[99]); 
    assign layer_0[7828] = ~in[583] | (in[452] & in[583]); 
    assign layer_0[7829] = ~in[295] | (in[295] & in[624]); 
    assign layer_0[7830] = ~in[35] | (in[229] & in[35]); 
    assign layer_0[7831] = ~in[480]; 
    assign layer_0[7832] = ~in[190] | (in[667] & in[190]); 
    assign layer_0[7833] = in[317] ^ in[488]; 
    assign layer_0[7834] = ~(in[204] ^ in[564]); 
    assign layer_0[7835] = ~(in[658] | in[492]); 
    assign layer_0[7836] = ~(in[490] | in[18]); 
    assign layer_0[7837] = in[85]; 
    assign layer_0[7838] = ~in[619] | (in[93] & in[619]); 
    assign layer_0[7839] = ~(in[544] | in[187]); 
    assign layer_0[7840] = in[339] ^ in[536]; 
    assign layer_0[7841] = in[29] ^ in[724]; 
    assign layer_0[7842] = ~in[682]; 
    assign layer_0[7843] = in[643] ^ in[205]; 
    assign layer_0[7844] = in[566] ^ in[453]; 
    assign layer_0[7845] = in[1] & ~in[7]; 
    assign layer_0[7846] = ~(in[472] ^ in[659]); 
    assign layer_0[7847] = ~in[612] | (in[722] & in[612]); 
    assign layer_0[7848] = ~(in[227] ^ in[706]); 
    assign layer_0[7849] = in[88]; 
    assign layer_0[7850] = ~(in[721] | in[504]); 
    assign layer_0[7851] = in[64] | in[420]; 
    assign layer_0[7852] = ~in[161]; 
    assign layer_0[7853] = in[236] | in[650]; 
    assign layer_0[7854] = ~(in[80] & in[347]); 
    assign layer_0[7855] = ~in[502] | (in[502] & in[501]); 
    assign layer_0[7856] = 1'b1; 
    assign layer_0[7857] = ~(in[315] ^ in[330]); 
    assign layer_0[7858] = ~in[603] | (in[62] & in[603]); 
    assign layer_0[7859] = ~in[679]; 
    assign layer_0[7860] = ~(in[558] ^ in[634]); 
    assign layer_0[7861] = ~(in[323] & in[65]); 
    assign layer_0[7862] = ~in[395] | (in[318] & in[395]); 
    assign layer_0[7863] = ~in[646] | (in[458] & in[646]); 
    assign layer_0[7864] = in[646] ^ in[647]; 
    assign layer_0[7865] = in[348] & in[650]; 
    assign layer_0[7866] = in[551] & ~in[634]; 
    assign layer_0[7867] = in[228] ^ in[246]; 
    assign layer_0[7868] = in[312] ^ in[692]; 
    assign layer_0[7869] = in[4] ^ in[53]; 
    assign layer_0[7870] = in[498] & ~in[527]; 
    assign layer_0[7871] = in[473] | in[645]; 
    assign layer_0[7872] = in[4] | in[671]; 
    assign layer_0[7873] = in[550] ^ in[565]; 
    assign layer_0[7874] = in[72]; 
    assign layer_0[7875] = ~(in[711] | in[712]); 
    assign layer_0[7876] = ~in[314] | (in[314] & in[657]); 
    assign layer_0[7877] = ~in[628] | (in[628] & in[588]); 
    assign layer_0[7878] = in[158] | in[491]; 
    assign layer_0[7879] = ~in[633]; 
    assign layer_0[7880] = in[190]; 
    assign layer_0[7881] = ~(in[246] ^ in[285]); 
    assign layer_0[7882] = in[715] | in[614]; 
    assign layer_0[7883] = ~(in[46] ^ in[18]); 
    assign layer_0[7884] = ~(in[662] & in[331]); 
    assign layer_0[7885] = ~(in[262] & in[18]); 
    assign layer_0[7886] = ~in[252]; 
    assign layer_0[7887] = in[308] & in[209]; 
    assign layer_0[7888] = ~(in[225] | in[47]); 
    assign layer_0[7889] = in[119] & in[249]; 
    assign layer_0[7890] = in[392]; 
    assign layer_0[7891] = in[508]; 
    assign layer_0[7892] = ~(in[761] ^ in[538]); 
    assign layer_0[7893] = in[728] & ~in[186]; 
    assign layer_0[7894] = in[280] & ~in[366]; 
    assign layer_0[7895] = in[506] ^ in[34]; 
    assign layer_0[7896] = in[580] ^ in[204]; 
    assign layer_0[7897] = ~(in[441] ^ in[264]); 
    assign layer_0[7898] = ~(in[322] ^ in[339]); 
    assign layer_0[7899] = in[709] ^ in[262]; 
    assign layer_0[7900] = ~(in[462] ^ in[488]); 
    assign layer_0[7901] = in[300] ^ in[597]; 
    assign layer_0[7902] = ~(in[180] & in[576]); 
    assign layer_0[7903] = in[61] ^ in[606]; 
    assign layer_0[7904] = in[599] ^ in[695]; 
    assign layer_0[7905] = ~(in[309] ^ in[487]); 
    assign layer_0[7906] = in[420] & ~in[505]; 
    assign layer_0[7907] = ~(in[710] & in[292]); 
    assign layer_0[7908] = in[84] ^ in[287]; 
    assign layer_0[7909] = ~(in[490] & in[121]); 
    assign layer_0[7910] = ~(in[622] ^ in[335]); 
    assign layer_0[7911] = ~in[598]; 
    assign layer_0[7912] = in[275]; 
    assign layer_0[7913] = in[523] ^ in[194]; 
    assign layer_0[7914] = in[341]; 
    assign layer_0[7915] = in[710] & ~in[174]; 
    assign layer_0[7916] = in[608] | in[742]; 
    assign layer_0[7917] = ~in[145] | (in[639] & in[145]); 
    assign layer_0[7918] = in[756] ^ in[215]; 
    assign layer_0[7919] = in[60] & in[123]; 
    assign layer_0[7920] = in[643] ^ in[651]; 
    assign layer_0[7921] = ~in[311] | (in[311] & in[173]); 
    assign layer_0[7922] = in[508] & in[296]; 
    assign layer_0[7923] = ~in[602] | (in[602] & in[620]); 
    assign layer_0[7924] = in[326]; 
    assign layer_0[7925] = in[438] & ~in[748]; 
    assign layer_0[7926] = in[325] & ~in[248]; 
    assign layer_0[7927] = ~(in[651] & in[281]); 
    assign layer_0[7928] = ~(in[50] & in[225]); 
    assign layer_0[7929] = in[472] & ~in[361]; 
    assign layer_0[7930] = ~in[62] | (in[70] & in[62]); 
    assign layer_0[7931] = ~(in[631] ^ in[632]); 
    assign layer_0[7932] = ~(in[373] | in[80]); 
    assign layer_0[7933] = in[310] ^ in[619]; 
    assign layer_0[7934] = ~(in[357] | in[371]); 
    assign layer_0[7935] = in[220] & in[401]; 
    assign layer_0[7936] = ~(in[482] ^ in[604]); 
    assign layer_0[7937] = ~in[570]; 
    assign layer_0[7938] = in[694] ^ in[695]; 
    assign layer_0[7939] = ~(in[111] ^ in[94]); 
    assign layer_0[7940] = in[230] & in[519]; 
    assign layer_0[7941] = ~in[3] | (in[3] & in[684]); 
    assign layer_0[7942] = ~(in[124] ^ in[580]); 
    assign layer_0[7943] = ~in[727] | (in[727] & in[386]); 
    assign layer_0[7944] = ~(in[629] ^ in[636]); 
    assign layer_0[7945] = in[331] ^ in[535]; 
    assign layer_0[7946] = in[348] & in[692]; 
    assign layer_0[7947] = in[398] & in[180]; 
    assign layer_0[7948] = ~in[5] | (in[452] & in[5]); 
    assign layer_0[7949] = in[507] | in[616]; 
    assign layer_0[7950] = ~in[566]; 
    assign layer_0[7951] = in[556] & ~in[674]; 
    assign layer_0[7952] = in[45] ^ in[281]; 
    assign layer_0[7953] = in[699]; 
    assign layer_0[7954] = ~(in[482] | in[175]); 
    assign layer_0[7955] = 1'b0; 
    assign layer_0[7956] = in[446] & ~in[757]; 
    assign layer_0[7957] = in[95] ^ in[24]; 
    assign layer_0[7958] = ~(in[98] | in[632]); 
    assign layer_0[7959] = ~(in[70] | in[114]); 
    assign layer_0[7960] = ~in[595]; 
    assign layer_0[7961] = ~(in[746] ^ in[612]); 
    assign layer_0[7962] = in[293]; 
    assign layer_0[7963] = in[28] ^ in[616]; 
    assign layer_0[7964] = ~in[252] | (in[461] & in[252]); 
    assign layer_0[7965] = in[185] | in[352]; 
    assign layer_0[7966] = ~(in[374] | in[587]); 
    assign layer_0[7967] = ~(in[276] & in[115]); 
    assign layer_0[7968] = in[628] ^ in[308]; 
    assign layer_0[7969] = ~in[724]; 
    assign layer_0[7970] = in[563]; 
    assign layer_0[7971] = ~in[329]; 
    assign layer_0[7972] = in[407] & ~in[575]; 
    assign layer_0[7973] = in[730] ^ in[33]; 
    assign layer_0[7974] = in[24] ^ in[319]; 
    assign layer_0[7975] = ~in[98]; 
    assign layer_0[7976] = ~(in[8] ^ in[156]); 
    assign layer_0[7977] = 1'b1; 
    assign layer_0[7978] = ~in[517] | (in[650] & in[517]); 
    assign layer_0[7979] = ~in[324] | (in[523] & in[324]); 
    assign layer_0[7980] = in[543]; 
    assign layer_0[7981] = in[85] & ~in[74]; 
    assign layer_0[7982] = ~in[264]; 
    assign layer_0[7983] = ~(in[762] ^ in[681]); 
    assign layer_0[7984] = in[280] | in[244]; 
    assign layer_0[7985] = in[732]; 
    assign layer_0[7986] = in[88] & ~in[672]; 
    assign layer_0[7987] = ~(in[751] ^ in[245]); 
    assign layer_0[7988] = in[40]; 
    assign layer_0[7989] = in[17] | in[536]; 
    assign layer_0[7990] = ~in[611]; 
    assign layer_0[7991] = ~(in[360] ^ in[344]); 
    assign layer_0[7992] = ~(in[694] | in[626]); 
    assign layer_0[7993] = ~(in[613] | in[516]); 
    assign layer_0[7994] = in[476] ^ in[4]; 
    assign layer_0[7995] = in[520] & ~in[137]; 
    assign layer_0[7996] = ~in[169]; 
    assign layer_0[7997] = in[586] ^ in[444]; 
    assign layer_0[7998] = in[324]; 
    assign layer_0[7999] = in[165] & in[11]; 
    // Layer 1 ============================================================
    assign out[0] = ~(layer_0[1967] ^ layer_0[2911]); 
    assign out[1] = layer_0[3120] | layer_0[7946]; 
    assign out[2] = ~(layer_0[7289] ^ layer_0[3989]); 
    assign out[3] = ~(layer_0[6853] ^ layer_0[506]); 
    assign out[4] = ~layer_0[1694]; 
    assign out[5] = layer_0[7638] & ~layer_0[4265]; 
    assign out[6] = layer_0[3523] ^ layer_0[3613]; 
    assign out[7] = layer_0[4310]; 
    assign out[8] = ~(layer_0[4400] ^ layer_0[2764]); 
    assign out[9] = ~(layer_0[2607] | layer_0[1513]); 
    assign out[10] = ~(layer_0[6754] & layer_0[2359]); 
    assign out[11] = layer_0[3495] | layer_0[1660]; 
    assign out[12] = layer_0[5205] & layer_0[7622]; 
    assign out[13] = ~(layer_0[6899] ^ layer_0[6487]); 
    assign out[14] = layer_0[195] | layer_0[5219]; 
    assign out[15] = ~layer_0[7864]; 
    assign out[16] = layer_0[4454] & ~layer_0[3498]; 
    assign out[17] = layer_0[4787]; 
    assign out[18] = ~(layer_0[5806] ^ layer_0[1558]); 
    assign out[19] = layer_0[5820] ^ layer_0[3722]; 
    assign out[20] = ~layer_0[1399] | (layer_0[2723] & layer_0[1399]); 
    assign out[21] = layer_0[6789]; 
    assign out[22] = layer_0[508] ^ layer_0[4131]; 
    assign out[23] = layer_0[4201] ^ layer_0[2066]; 
    assign out[24] = layer_0[7057] ^ layer_0[7524]; 
    assign out[25] = ~(layer_0[4158] & layer_0[2333]); 
    assign out[26] = ~layer_0[4322]; 
    assign out[27] = ~(layer_0[785] ^ layer_0[2163]); 
    assign out[28] = layer_0[190]; 
    assign out[29] = layer_0[3507] ^ layer_0[183]; 
    assign out[30] = layer_0[1169] ^ layer_0[5979]; 
    assign out[31] = layer_0[7454] & ~layer_0[7069]; 
    assign out[32] = layer_0[5830] ^ layer_0[6902]; 
    assign out[33] = ~layer_0[4875]; 
    assign out[34] = layer_0[2783] ^ layer_0[6303]; 
    assign out[35] = layer_0[2647]; 
    assign out[36] = layer_0[2345] & layer_0[2015]; 
    assign out[37] = layer_0[7113] ^ layer_0[4215]; 
    assign out[38] = ~layer_0[2612]; 
    assign out[39] = ~(layer_0[608] & layer_0[7257]); 
    assign out[40] = ~(layer_0[3234] ^ layer_0[262]); 
    assign out[41] = layer_0[3005]; 
    assign out[42] = layer_0[3361] ^ layer_0[5646]; 
    assign out[43] = ~(layer_0[1445] | layer_0[4461]); 
    assign out[44] = ~layer_0[4089]; 
    assign out[45] = layer_0[5141] ^ layer_0[238]; 
    assign out[46] = layer_0[5001] ^ layer_0[856]; 
    assign out[47] = layer_0[4651] ^ layer_0[5258]; 
    assign out[48] = ~(layer_0[1215] & layer_0[7716]); 
    assign out[49] = ~(layer_0[626] & layer_0[466]); 
    assign out[50] = layer_0[6391] ^ layer_0[2048]; 
    assign out[51] = ~(layer_0[3790] ^ layer_0[7936]); 
    assign out[52] = layer_0[4368] | layer_0[3253]; 
    assign out[53] = ~(layer_0[4904] ^ layer_0[1653]); 
    assign out[54] = layer_0[5084] | layer_0[5168]; 
    assign out[55] = layer_0[5720] & ~layer_0[4159]; 
    assign out[56] = ~(layer_0[5788] ^ layer_0[4775]); 
    assign out[57] = layer_0[3394] & ~layer_0[168]; 
    assign out[58] = ~layer_0[29] | (layer_0[1568] & layer_0[29]); 
    assign out[59] = ~(layer_0[1509] ^ layer_0[3224]); 
    assign out[60] = layer_0[3704] & ~layer_0[7744]; 
    assign out[61] = layer_0[3633]; 
    assign out[62] = layer_0[4177]; 
    assign out[63] = ~(layer_0[4263] & layer_0[3670]); 
    assign out[64] = ~layer_0[1323]; 
    assign out[65] = ~(layer_0[7779] ^ layer_0[4400]); 
    assign out[66] = ~layer_0[4539]; 
    assign out[67] = layer_0[7809] | layer_0[1711]; 
    assign out[68] = ~(layer_0[500] ^ layer_0[1034]); 
    assign out[69] = layer_0[7500] ^ layer_0[7961]; 
    assign out[70] = ~layer_0[4949] | (layer_0[6828] & layer_0[4949]); 
    assign out[71] = layer_0[4470] ^ layer_0[5209]; 
    assign out[72] = ~(layer_0[4016] ^ layer_0[7647]); 
    assign out[73] = ~layer_0[4074] | (layer_0[4074] & layer_0[4727]); 
    assign out[74] = layer_0[319] ^ layer_0[1726]; 
    assign out[75] = ~(layer_0[6855] ^ layer_0[6555]); 
    assign out[76] = layer_0[7662] ^ layer_0[5849]; 
    assign out[77] = ~(layer_0[2566] ^ layer_0[7274]); 
    assign out[78] = ~layer_0[1493]; 
    assign out[79] = layer_0[2377] ^ layer_0[6887]; 
    assign out[80] = layer_0[6821] | layer_0[5885]; 
    assign out[81] = ~layer_0[1379] | (layer_0[7115] & layer_0[1379]); 
    assign out[82] = layer_0[5619] ^ layer_0[910]; 
    assign out[83] = layer_0[4871] & ~layer_0[942]; 
    assign out[84] = layer_0[4161] | layer_0[6846]; 
    assign out[85] = layer_0[5603] & ~layer_0[3334]; 
    assign out[86] = layer_0[1491] & ~layer_0[1719]; 
    assign out[87] = ~layer_0[6199]; 
    assign out[88] = layer_0[5399] & layer_0[5465]; 
    assign out[89] = ~(layer_0[3196] ^ layer_0[5260]); 
    assign out[90] = ~(layer_0[4340] ^ layer_0[5297]); 
    assign out[91] = ~(layer_0[1968] ^ layer_0[5695]); 
    assign out[92] = ~layer_0[3460]; 
    assign out[93] = layer_0[5964] ^ layer_0[4420]; 
    assign out[94] = ~(layer_0[3126] ^ layer_0[7275]); 
    assign out[95] = layer_0[3150] ^ layer_0[3519]; 
    assign out[96] = ~layer_0[7461]; 
    assign out[97] = layer_0[6951] ^ layer_0[4062]; 
    assign out[98] = ~layer_0[7541]; 
    assign out[99] = layer_0[7223] ^ layer_0[4644]; 
    assign out[100] = ~(layer_0[7346] | layer_0[3565]); 
    assign out[101] = layer_0[3664] & layer_0[1199]; 
    assign out[102] = ~(layer_0[6576] & layer_0[3786]); 
    assign out[103] = ~layer_0[4195] | (layer_0[4195] & layer_0[1268]); 
    assign out[104] = ~(layer_0[4500] ^ layer_0[4969]); 
    assign out[105] = ~(layer_0[5281] ^ layer_0[266]); 
    assign out[106] = layer_0[4090] ^ layer_0[7260]; 
    assign out[107] = layer_0[1674] ^ layer_0[4306]; 
    assign out[108] = ~(layer_0[2491] ^ layer_0[7137]); 
    assign out[109] = layer_0[7425] ^ layer_0[7052]; 
    assign out[110] = layer_0[1421] ^ layer_0[5093]; 
    assign out[111] = ~layer_0[6489]; 
    assign out[112] = layer_0[1525] & ~layer_0[7302]; 
    assign out[113] = layer_0[2582] | layer_0[4671]; 
    assign out[114] = ~layer_0[5079] | (layer_0[3220] & layer_0[5079]); 
    assign out[115] = layer_0[4872]; 
    assign out[116] = layer_0[715] ^ layer_0[946]; 
    assign out[117] = ~(layer_0[3760] & layer_0[3644]); 
    assign out[118] = ~(layer_0[3506] ^ layer_0[5666]); 
    assign out[119] = ~(layer_0[7324] ^ layer_0[471]); 
    assign out[120] = layer_0[4900] ^ layer_0[5051]; 
    assign out[121] = ~layer_0[4071] | (layer_0[3346] & layer_0[4071]); 
    assign out[122] = ~(layer_0[1028] ^ layer_0[7997]); 
    assign out[123] = ~(layer_0[7338] ^ layer_0[6658]); 
    assign out[124] = ~layer_0[5019]; 
    assign out[125] = layer_0[6844] ^ layer_0[2559]; 
    assign out[126] = ~layer_0[1657] | (layer_0[1657] & layer_0[7310]); 
    assign out[127] = ~(layer_0[6917] ^ layer_0[2425]); 
    assign out[128] = layer_0[4199] & ~layer_0[668]; 
    assign out[129] = ~(layer_0[9] ^ layer_0[4097]); 
    assign out[130] = ~(layer_0[3399] ^ layer_0[7149]); 
    assign out[131] = ~(layer_0[3729] | layer_0[1091]); 
    assign out[132] = ~layer_0[6614]; 
    assign out[133] = ~(layer_0[1387] | layer_0[5829]); 
    assign out[134] = layer_0[6830] ^ layer_0[4219]; 
    assign out[135] = ~(layer_0[1598] ^ layer_0[4049]); 
    assign out[136] = layer_0[2696] ^ layer_0[518]; 
    assign out[137] = ~(layer_0[2141] ^ layer_0[5133]); 
    assign out[138] = ~(layer_0[4896] ^ layer_0[3512]); 
    assign out[139] = ~(layer_0[3163] ^ layer_0[4208]); 
    assign out[140] = ~layer_0[5984] | (layer_0[5984] & layer_0[2149]); 
    assign out[141] = ~(layer_0[2968] | layer_0[2330]); 
    assign out[142] = layer_0[6781] | layer_0[807]; 
    assign out[143] = layer_0[571] ^ layer_0[7302]; 
    assign out[144] = layer_0[5713] | layer_0[176]; 
    assign out[145] = layer_0[6474] ^ layer_0[7794]; 
    assign out[146] = layer_0[1727] ^ layer_0[6861]; 
    assign out[147] = ~layer_0[5158]; 
    assign out[148] = ~(layer_0[1472] ^ layer_0[3272]); 
    assign out[149] = ~(layer_0[3096] ^ layer_0[7331]); 
    assign out[150] = layer_0[894] | layer_0[602]; 
    assign out[151] = ~layer_0[516] | (layer_0[2285] & layer_0[516]); 
    assign out[152] = layer_0[1631] ^ layer_0[1009]; 
    assign out[153] = ~layer_0[1004]; 
    assign out[154] = layer_0[4540] & ~layer_0[4377]; 
    assign out[155] = layer_0[3378] ^ layer_0[3833]; 
    assign out[156] = layer_0[1626]; 
    assign out[157] = layer_0[7388] & ~layer_0[4905]; 
    assign out[158] = layer_0[3431] & ~layer_0[4480]; 
    assign out[159] = ~(layer_0[3614] | layer_0[2397]); 
    assign out[160] = ~(layer_0[2234] & layer_0[7698]); 
    assign out[161] = ~(layer_0[100] ^ layer_0[7506]); 
    assign out[162] = ~layer_0[7969] | (layer_0[5838] & layer_0[7969]); 
    assign out[163] = layer_0[7741]; 
    assign out[164] = layer_0[6952] & layer_0[4138]; 
    assign out[165] = ~(layer_0[94] ^ layer_0[1402]); 
    assign out[166] = layer_0[3858] ^ layer_0[884]; 
    assign out[167] = ~(layer_0[4136] ^ layer_0[4549]); 
    assign out[168] = layer_0[7721] ^ layer_0[1030]; 
    assign out[169] = layer_0[4435] ^ layer_0[3558]; 
    assign out[170] = ~layer_0[1219]; 
    assign out[171] = layer_0[909] ^ layer_0[5515]; 
    assign out[172] = layer_0[7491] & ~layer_0[6104]; 
    assign out[173] = layer_0[4650] ^ layer_0[2965]; 
    assign out[174] = layer_0[6773] ^ layer_0[1495]; 
    assign out[175] = layer_0[2235] ^ layer_0[464]; 
    assign out[176] = layer_0[4313] ^ layer_0[1618]; 
    assign out[177] = ~(layer_0[556] | layer_0[3089]); 
    assign out[178] = layer_0[2003] ^ layer_0[6557]; 
    assign out[179] = layer_0[342] ^ layer_0[3576]; 
    assign out[180] = ~layer_0[7870] | (layer_0[308] & layer_0[7870]); 
    assign out[181] = ~layer_0[3434]; 
    assign out[182] = ~(layer_0[7048] | layer_0[2278]); 
    assign out[183] = ~layer_0[3274] | (layer_0[3274] & layer_0[1594]); 
    assign out[184] = layer_0[7253]; 
    assign out[185] = ~layer_0[5994]; 
    assign out[186] = ~(layer_0[7694] ^ layer_0[5004]); 
    assign out[187] = layer_0[2413] ^ layer_0[5315]; 
    assign out[188] = ~(layer_0[4040] | layer_0[7763]); 
    assign out[189] = layer_0[2973] & ~layer_0[5663]; 
    assign out[190] = ~(layer_0[7963] ^ layer_0[743]); 
    assign out[191] = layer_0[4287] & ~layer_0[7834]; 
    assign out[192] = layer_0[2093] & ~layer_0[5953]; 
    assign out[193] = layer_0[2916] ^ layer_0[2531]; 
    assign out[194] = layer_0[6050] ^ layer_0[1894]; 
    assign out[195] = layer_0[6541]; 
    assign out[196] = layer_0[7173] & ~layer_0[2023]; 
    assign out[197] = ~layer_0[6239]; 
    assign out[198] = ~layer_0[1133]; 
    assign out[199] = ~(layer_0[5684] & layer_0[5]); 
    assign out[200] = ~(layer_0[3174] | layer_0[6689]); 
    assign out[201] = layer_0[4814] ^ layer_0[6017]; 
    assign out[202] = layer_0[6287] & layer_0[110]; 
    assign out[203] = ~(layer_0[4072] | layer_0[6799]); 
    assign out[204] = layer_0[4677] ^ layer_0[1015]; 
    assign out[205] = layer_0[3020] & ~layer_0[4192]; 
    assign out[206] = layer_0[1038] & ~layer_0[6383]; 
    assign out[207] = ~(layer_0[7932] | layer_0[5250]); 
    assign out[208] = layer_0[2864] & ~layer_0[5652]; 
    assign out[209] = ~layer_0[6775]; 
    assign out[210] = layer_0[7068] & ~layer_0[412]; 
    assign out[211] = layer_0[7913] ^ layer_0[1632]; 
    assign out[212] = layer_0[63] ^ layer_0[708]; 
    assign out[213] = layer_0[4190] & ~layer_0[2926]; 
    assign out[214] = ~(layer_0[4476] ^ layer_0[4399]); 
    assign out[215] = ~(layer_0[2961] ^ layer_0[4579]); 
    assign out[216] = layer_0[2310] ^ layer_0[5527]; 
    assign out[217] = layer_0[7968] ^ layer_0[1007]; 
    assign out[218] = ~(layer_0[2960] | layer_0[692]); 
    assign out[219] = layer_0[5584] ^ layer_0[4174]; 
    assign out[220] = layer_0[5480] & ~layer_0[4695]; 
    assign out[221] = layer_0[4682] ^ layer_0[4772]; 
    assign out[222] = layer_0[7083] ^ layer_0[5058]; 
    assign out[223] = layer_0[6231] ^ layer_0[4879]; 
    assign out[224] = layer_0[1354] & ~layer_0[3502]; 
    assign out[225] = ~(layer_0[4485] ^ layer_0[7067]); 
    assign out[226] = layer_0[1065] ^ layer_0[3047]; 
    assign out[227] = ~layer_0[6067]; 
    assign out[228] = layer_0[3703]; 
    assign out[229] = layer_0[1515]; 
    assign out[230] = ~(layer_0[173] ^ layer_0[4397]); 
    assign out[231] = layer_0[6699] ^ layer_0[5532]; 
    assign out[232] = layer_0[259] ^ layer_0[1400]; 
    assign out[233] = ~(layer_0[6503] | layer_0[3315]); 
    assign out[234] = layer_0[1291] & ~layer_0[4559]; 
    assign out[235] = ~(layer_0[701] ^ layer_0[6992]); 
    assign out[236] = ~layer_0[3429] | (layer_0[3429] & layer_0[92]); 
    assign out[237] = ~layer_0[5082] | (layer_0[476] & layer_0[5082]); 
    assign out[238] = layer_0[4370] | layer_0[7227]; 
    assign out[239] = layer_0[5022]; 
    assign out[240] = ~(layer_0[7942] ^ layer_0[7574]); 
    assign out[241] = ~layer_0[5785] | (layer_0[1254] & layer_0[5785]); 
    assign out[242] = layer_0[7620] ^ layer_0[4321]; 
    assign out[243] = ~layer_0[2746] | (layer_0[2746] & layer_0[4933]); 
    assign out[244] = ~layer_0[6857] | (layer_0[6857] & layer_0[2376]); 
    assign out[245] = ~(layer_0[3283] ^ layer_0[7071]); 
    assign out[246] = ~(layer_0[5819] ^ layer_0[5947]); 
    assign out[247] = layer_0[5965] ^ layer_0[2240]; 
    assign out[248] = layer_0[6544] ^ layer_0[3685]; 
    assign out[249] = ~layer_0[848] | (layer_0[848] & layer_0[2052]); 
    assign out[250] = layer_0[339] | layer_0[5575]; 
    assign out[251] = ~layer_0[3658] | (layer_0[7680] & layer_0[3658]); 
    assign out[252] = ~(layer_0[6493] ^ layer_0[7927]); 
    assign out[253] = ~layer_0[6009]; 
    assign out[254] = ~(layer_0[4998] ^ layer_0[7355]); 
    assign out[255] = layer_0[2364] ^ layer_0[2702]; 
    assign out[256] = layer_0[6794] ^ layer_0[5025]; 
    assign out[257] = ~(layer_0[4864] ^ layer_0[2378]); 
    assign out[258] = ~layer_0[3909]; 
    assign out[259] = ~(layer_0[6691] ^ layer_0[7511]); 
    assign out[260] = ~(layer_0[6895] ^ layer_0[1705]); 
    assign out[261] = ~(layer_0[844] ^ layer_0[638]); 
    assign out[262] = layer_0[804] | layer_0[6561]; 
    assign out[263] = layer_0[6154] ^ layer_0[1707]; 
    assign out[264] = layer_0[2732] ^ layer_0[1781]; 
    assign out[265] = ~(layer_0[4652] ^ layer_0[2162]); 
    assign out[266] = ~layer_0[16] | (layer_0[1482] & layer_0[16]); 
    assign out[267] = ~(layer_0[7086] ^ layer_0[126]); 
    assign out[268] = layer_0[170] ^ layer_0[4171]; 
    assign out[269] = ~(layer_0[1990] ^ layer_0[3107]); 
    assign out[270] = layer_0[3995] ^ layer_0[3545]; 
    assign out[271] = ~(layer_0[6540] & layer_0[955]); 
    assign out[272] = ~layer_0[411] | (layer_0[7039] & layer_0[411]); 
    assign out[273] = layer_0[3084] ^ layer_0[68]; 
    assign out[274] = ~layer_0[2248] | (layer_0[2248] & layer_0[3397]); 
    assign out[275] = layer_0[898] ^ layer_0[3353]; 
    assign out[276] = ~layer_0[1845] | (layer_0[5930] & layer_0[1845]); 
    assign out[277] = layer_0[3233] ^ layer_0[4212]; 
    assign out[278] = ~(layer_0[5014] ^ layer_0[7487]); 
    assign out[279] = layer_0[2291]; 
    assign out[280] = ~(layer_0[3969] ^ layer_0[2841]); 
    assign out[281] = layer_0[6319]; 
    assign out[282] = layer_0[3887]; 
    assign out[283] = ~(layer_0[1039] ^ layer_0[1736]); 
    assign out[284] = ~(layer_0[3050] ^ layer_0[7658]); 
    assign out[285] = layer_0[1251] ^ layer_0[2215]; 
    assign out[286] = layer_0[4041] | layer_0[4311]; 
    assign out[287] = ~(layer_0[7686] ^ layer_0[7659]); 
    assign out[288] = layer_0[2119]; 
    assign out[289] = layer_0[5385] | layer_0[7247]; 
    assign out[290] = ~(layer_0[2252] ^ layer_0[2852]); 
    assign out[291] = layer_0[3325] & layer_0[1761]; 
    assign out[292] = ~(layer_0[1489] ^ layer_0[6858]); 
    assign out[293] = ~layer_0[7607]; 
    assign out[294] = layer_0[5916] ^ layer_0[6227]; 
    assign out[295] = layer_0[1262]; 
    assign out[296] = layer_0[4971]; 
    assign out[297] = ~(layer_0[1081] ^ layer_0[1404]); 
    assign out[298] = layer_0[1330] ^ layer_0[5774]; 
    assign out[299] = layer_0[2819]; 
    assign out[300] = layer_0[3625]; 
    assign out[301] = layer_0[6367]; 
    assign out[302] = layer_0[3748] ^ layer_0[7963]; 
    assign out[303] = layer_0[5959] ^ layer_0[2966]; 
    assign out[304] = ~(layer_0[5427] & layer_0[4037]); 
    assign out[305] = ~layer_0[7190]; 
    assign out[306] = layer_0[248] ^ layer_0[7784]; 
    assign out[307] = layer_0[6709] ^ layer_0[2501]; 
    assign out[308] = layer_0[5542] & ~layer_0[6074]; 
    assign out[309] = layer_0[6148] & layer_0[1988]; 
    assign out[310] = layer_0[6798]; 
    assign out[311] = layer_0[4809] ^ layer_0[2449]; 
    assign out[312] = layer_0[2845] & ~layer_0[4718]; 
    assign out[313] = ~(layer_0[3686] ^ layer_0[5544]); 
    assign out[314] = ~layer_0[6713] | (layer_0[6713] & layer_0[7906]); 
    assign out[315] = layer_0[2592] & layer_0[7358]; 
    assign out[316] = ~layer_0[5007] | (layer_0[3745] & layer_0[5007]); 
    assign out[317] = layer_0[5382] ^ layer_0[4002]; 
    assign out[318] = layer_0[7628] ^ layer_0[5053]; 
    assign out[319] = ~(layer_0[413] ^ layer_0[5690]); 
    assign out[320] = layer_0[4979] ^ layer_0[1141]; 
    assign out[321] = layer_0[6808] | layer_0[2528]; 
    assign out[322] = layer_0[2379] ^ layer_0[3295]; 
    assign out[323] = layer_0[7055]; 
    assign out[324] = layer_0[1580] ^ layer_0[4039]; 
    assign out[325] = layer_0[3145] | layer_0[3480]; 
    assign out[326] = ~(layer_0[6921] ^ layer_0[3373]); 
    assign out[327] = ~(layer_0[7748] & layer_0[5871]); 
    assign out[328] = layer_0[846] & layer_0[7529]; 
    assign out[329] = ~layer_0[2677] | (layer_0[2677] & layer_0[3010]); 
    assign out[330] = ~(layer_0[1411] ^ layer_0[1472]); 
    assign out[331] = ~(layer_0[522] ^ layer_0[5578]); 
    assign out[332] = layer_0[7661] & ~layer_0[1342]; 
    assign out[333] = layer_0[5337]; 
    assign out[334] = layer_0[5839] ^ layer_0[2544]; 
    assign out[335] = layer_0[6212] ^ layer_0[1048]; 
    assign out[336] = layer_0[6128] ^ layer_0[4567]; 
    assign out[337] = layer_0[4121] ^ layer_0[3117]; 
    assign out[338] = ~(layer_0[1859] | layer_0[4039]); 
    assign out[339] = ~layer_0[5702] | (layer_0[5702] & layer_0[5667]); 
    assign out[340] = ~(layer_0[7879] ^ layer_0[2440]); 
    assign out[341] = ~(layer_0[6458] ^ layer_0[3575]); 
    assign out[342] = layer_0[6025] ^ layer_0[5855]; 
    assign out[343] = layer_0[2288] ^ layer_0[5856]; 
    assign out[344] = ~(layer_0[5563] | layer_0[7091]); 
    assign out[345] = ~layer_0[257] | (layer_0[7248] & layer_0[257]); 
    assign out[346] = layer_0[6937] ^ layer_0[1002]; 
    assign out[347] = ~(layer_0[5722] ^ layer_0[3113]); 
    assign out[348] = layer_0[3077]; 
    assign out[349] = ~(layer_0[5710] ^ layer_0[6421]); 
    assign out[350] = layer_0[6827]; 
    assign out[351] = layer_0[7383]; 
    assign out[352] = layer_0[3205] ^ layer_0[5354]; 
    assign out[353] = layer_0[5128] & ~layer_0[2118]; 
    assign out[354] = ~(layer_0[2368] ^ layer_0[711]); 
    assign out[355] = layer_0[5319] & ~layer_0[3339]; 
    assign out[356] = layer_0[2596] & ~layer_0[6317]; 
    assign out[357] = layer_0[202] & ~layer_0[5741]; 
    assign out[358] = ~layer_0[5378]; 
    assign out[359] = ~layer_0[4639] | (layer_0[4639] & layer_0[4894]); 
    assign out[360] = layer_0[259] | layer_0[6789]; 
    assign out[361] = ~(layer_0[1315] | layer_0[6021]); 
    assign out[362] = layer_0[3718] & ~layer_0[1146]; 
    assign out[363] = ~layer_0[7866] | (layer_0[7866] & layer_0[1922]); 
    assign out[364] = layer_0[3926] ^ layer_0[1087]; 
    assign out[365] = layer_0[2058]; 
    assign out[366] = layer_0[13]; 
    assign out[367] = layer_0[4034] ^ layer_0[7663]; 
    assign out[368] = layer_0[1722]; 
    assign out[369] = layer_0[5902] | layer_0[4253]; 
    assign out[370] = ~layer_0[4007] | (layer_0[658] & layer_0[4007]); 
    assign out[371] = layer_0[5109]; 
    assign out[372] = layer_0[7825] ^ layer_0[7448]; 
    assign out[373] = ~layer_0[5208]; 
    assign out[374] = layer_0[5675]; 
    assign out[375] = layer_0[7510] ^ layer_0[5501]; 
    assign out[376] = layer_0[3792] ^ layer_0[6375]; 
    assign out[377] = ~(layer_0[7143] ^ layer_0[1346]); 
    assign out[378] = ~layer_0[385] | (layer_0[1991] & layer_0[385]); 
    assign out[379] = ~layer_0[488]; 
    assign out[380] = layer_0[293] & layer_0[5247]; 
    assign out[381] = layer_0[1463] ^ layer_0[4665]; 
    assign out[382] = layer_0[7177] ^ layer_0[4284]; 
    assign out[383] = ~(layer_0[903] ^ layer_0[7742]); 
    assign out[384] = ~(layer_0[6746] & layer_0[5300]); 
    assign out[385] = layer_0[2306] ^ layer_0[366]; 
    assign out[386] = layer_0[4609] & layer_0[7514]; 
    assign out[387] = ~(layer_0[323] ^ layer_0[1134]); 
    assign out[388] = ~(layer_0[1826] & layer_0[6062]); 
    assign out[389] = layer_0[7319] ^ layer_0[3724]; 
    assign out[390] = layer_0[7692] | layer_0[5335]; 
    assign out[391] = ~layer_0[341] | (layer_0[341] & layer_0[1798]); 
    assign out[392] = layer_0[5162] ^ layer_0[7386]; 
    assign out[393] = layer_0[7370] ^ layer_0[1192]; 
    assign out[394] = layer_0[2465] & ~layer_0[5277]; 
    assign out[395] = ~layer_0[4997]; 
    assign out[396] = layer_0[225] ^ layer_0[6883]; 
    assign out[397] = layer_0[3369] ^ layer_0[7846]; 
    assign out[398] = layer_0[1459] ^ layer_0[1276]; 
    assign out[399] = ~(layer_0[953] | layer_0[3074]); 
    assign out[400] = layer_0[5921] | layer_0[1646]; 
    assign out[401] = layer_0[7640] ^ layer_0[7219]; 
    assign out[402] = ~(layer_0[5782] ^ layer_0[7153]); 
    assign out[403] = layer_0[5238] ^ layer_0[916]; 
    assign out[404] = ~(layer_0[6917] | layer_0[6593]); 
    assign out[405] = ~(layer_0[5835] ^ layer_0[1607]); 
    assign out[406] = layer_0[1436] & layer_0[2922]; 
    assign out[407] = ~layer_0[1878] | (layer_0[584] & layer_0[1878]); 
    assign out[408] = layer_0[3191] ^ layer_0[4385]; 
    assign out[409] = ~layer_0[2728] | (layer_0[2728] & layer_0[7463]); 
    assign out[410] = layer_0[5561] ^ layer_0[354]; 
    assign out[411] = ~(layer_0[1089] ^ layer_0[1076]); 
    assign out[412] = ~(layer_0[3738] | layer_0[902]); 
    assign out[413] = ~(layer_0[7820] ^ layer_0[6796]); 
    assign out[414] = ~(layer_0[4422] | layer_0[4844]); 
    assign out[415] = ~(layer_0[1739] ^ layer_0[7053]); 
    assign out[416] = layer_0[1564] ^ layer_0[6439]; 
    assign out[417] = layer_0[1695]; 
    assign out[418] = layer_0[6726]; 
    assign out[419] = layer_0[4112] & layer_0[749]; 
    assign out[420] = ~(layer_0[4897] ^ layer_0[292]); 
    assign out[421] = layer_0[7814] ^ layer_0[7954]; 
    assign out[422] = layer_0[5733] ^ layer_0[3448]; 
    assign out[423] = ~(layer_0[5112] ^ layer_0[2931]); 
    assign out[424] = 1'b1; 
    assign out[425] = ~layer_0[4167]; 
    assign out[426] = layer_0[2137]; 
    assign out[427] = layer_0[5138]; 
    assign out[428] = ~(layer_0[644] ^ layer_0[5605]); 
    assign out[429] = ~layer_0[7111]; 
    assign out[430] = ~layer_0[144] | (layer_0[144] & layer_0[7751]); 
    assign out[431] = ~(layer_0[4598] ^ layer_0[2210]); 
    assign out[432] = layer_0[6662] ^ layer_0[4254]; 
    assign out[433] = ~(layer_0[4592] & layer_0[1621]); 
    assign out[434] = ~(layer_0[2862] ^ layer_0[4141]); 
    assign out[435] = layer_0[5587] & ~layer_0[5671]; 
    assign out[436] = layer_0[7639] | layer_0[4163]; 
    assign out[437] = layer_0[4937] | layer_0[5188]; 
    assign out[438] = ~(layer_0[3868] ^ layer_0[7644]); 
    assign out[439] = ~(layer_0[6004] ^ layer_0[5911]); 
    assign out[440] = layer_0[1322] ^ layer_0[3637]; 
    assign out[441] = layer_0[1351] | layer_0[1366]; 
    assign out[442] = ~(layer_0[6605] ^ layer_0[326]); 
    assign out[443] = layer_0[6819] ^ layer_0[5143]; 
    assign out[444] = layer_0[1714] & ~layer_0[680]; 
    assign out[445] = layer_0[4820] ^ layer_0[1640]; 
    assign out[446] = ~(layer_0[5976] ^ layer_0[2967]); 
    assign out[447] = layer_0[371] ^ layer_0[6411]; 
    assign out[448] = ~(layer_0[7941] ^ layer_0[5376]); 
    assign out[449] = ~(layer_0[1607] ^ layer_0[2134]); 
    assign out[450] = layer_0[7084] ^ layer_0[4568]; 
    assign out[451] = ~(layer_0[662] ^ layer_0[1056]); 
    assign out[452] = layer_0[6121] ^ layer_0[7146]; 
    assign out[453] = layer_0[7899] ^ layer_0[7836]; 
    assign out[454] = ~(layer_0[5469] & layer_0[4799]); 
    assign out[455] = ~layer_0[4185] | (layer_0[5087] & layer_0[4185]); 
    assign out[456] = layer_0[5769] & layer_0[2504]; 
    assign out[457] = ~(layer_0[399] ^ layer_0[857]); 
    assign out[458] = ~(layer_0[6635] ^ layer_0[1499]); 
    assign out[459] = ~layer_0[4826]; 
    assign out[460] = ~(layer_0[7662] & layer_0[3867]); 
    assign out[461] = layer_0[1940] ^ layer_0[3608]; 
    assign out[462] = layer_0[2743] ^ layer_0[3607]; 
    assign out[463] = layer_0[4576] ^ layer_0[7206]; 
    assign out[464] = layer_0[6910] ^ layer_0[1548]; 
    assign out[465] = layer_0[5557]; 
    assign out[466] = ~layer_0[4053] | (layer_0[4964] & layer_0[4053]); 
    assign out[467] = ~(layer_0[2709] ^ layer_0[4186]); 
    assign out[468] = ~layer_0[1324]; 
    assign out[469] = ~(layer_0[2191] ^ layer_0[4685]); 
    assign out[470] = layer_0[4719] & layer_0[1954]; 
    assign out[471] = ~(layer_0[6431] | layer_0[1844]); 
    assign out[472] = ~(layer_0[6990] ^ layer_0[5761]); 
    assign out[473] = layer_0[507] & layer_0[231]; 
    assign out[474] = layer_0[7004] & ~layer_0[1741]; 
    assign out[475] = layer_0[156] & ~layer_0[6886]; 
    assign out[476] = layer_0[6485] ^ layer_0[6717]; 
    assign out[477] = ~(layer_0[1303] ^ layer_0[5789]); 
    assign out[478] = layer_0[4787]; 
    assign out[479] = ~layer_0[1816]; 
    assign out[480] = ~(layer_0[5478] & layer_0[2150]); 
    assign out[481] = ~(layer_0[5404] ^ layer_0[7698]); 
    assign out[482] = layer_0[1061] ^ layer_0[881]; 
    assign out[483] = ~(layer_0[266] ^ layer_0[7096]); 
    assign out[484] = layer_0[1523] & ~layer_0[340]; 
    assign out[485] = ~(layer_0[2035] ^ layer_0[6734]); 
    assign out[486] = ~(layer_0[7843] ^ layer_0[7311]); 
    assign out[487] = ~(layer_0[2176] ^ layer_0[6571]); 
    assign out[488] = layer_0[6731] & layer_0[7648]; 
    assign out[489] = ~layer_0[1583] | (layer_0[1583] & layer_0[6949]); 
    assign out[490] = layer_0[3385] | layer_0[7944]; 
    assign out[491] = layer_0[6301]; 
    assign out[492] = layer_0[3106] ^ layer_0[6157]; 
    assign out[493] = ~(layer_0[5181] & layer_0[2638]); 
    assign out[494] = ~layer_0[1673] | (layer_0[5318] & layer_0[1673]); 
    assign out[495] = ~(layer_0[1336] ^ layer_0[2722]); 
    assign out[496] = ~(layer_0[4705] ^ layer_0[6855]); 
    assign out[497] = layer_0[4989] ^ layer_0[1964]; 
    assign out[498] = ~layer_0[3592]; 
    assign out[499] = layer_0[2021]; 
    assign out[500] = ~layer_0[2017]; 
    assign out[501] = layer_0[1108] ^ layer_0[959]; 
    assign out[502] = layer_0[3263] | layer_0[7604]; 
    assign out[503] = layer_0[6940] & layer_0[3542]; 
    assign out[504] = layer_0[4634] ^ layer_0[2932]; 
    assign out[505] = layer_0[7132] ^ layer_0[6963]; 
    assign out[506] = ~(layer_0[6995] | layer_0[7367]); 
    assign out[507] = layer_0[6335] ^ layer_0[5744]; 
    assign out[508] = layer_0[845] | layer_0[4830]; 
    assign out[509] = layer_0[6873] ^ layer_0[253]; 
    assign out[510] = layer_0[2604] | layer_0[1405]; 
    assign out[511] = ~(layer_0[5391] ^ layer_0[7109]); 
    assign out[512] = ~(layer_0[3688] ^ layer_0[7046]); 
    assign out[513] = ~(layer_0[7509] ^ layer_0[317]); 
    assign out[514] = ~layer_0[4524] | (layer_0[7708] & layer_0[4524]); 
    assign out[515] = ~layer_0[6675]; 
    assign out[516] = layer_0[4999] ^ layer_0[2318]; 
    assign out[517] = ~layer_0[3363]; 
    assign out[518] = layer_0[1806] ^ layer_0[4860]; 
    assign out[519] = layer_0[1956] & ~layer_0[4819]; 
    assign out[520] = layer_0[1086] & ~layer_0[1494]; 
    assign out[521] = ~layer_0[1569] | (layer_0[1569] & layer_0[2626]); 
    assign out[522] = layer_0[5740] ^ layer_0[5750]; 
    assign out[523] = layer_0[5847] & layer_0[6604]; 
    assign out[524] = ~layer_0[1723] | (layer_0[5415] & layer_0[1723]); 
    assign out[525] = ~layer_0[6911]; 
    assign out[526] = layer_0[6357] & layer_0[215]; 
    assign out[527] = ~(layer_0[7207] ^ layer_0[7387]); 
    assign out[528] = layer_0[96] ^ layer_0[7612]; 
    assign out[529] = layer_0[7384] & ~layer_0[6968]; 
    assign out[530] = layer_0[3124] & ~layer_0[1017]; 
    assign out[531] = ~(layer_0[3273] & layer_0[6495]); 
    assign out[532] = ~(layer_0[5629] ^ layer_0[2498]); 
    assign out[533] = layer_0[5680]; 
    assign out[534] = layer_0[2497] & ~layer_0[2557]; 
    assign out[535] = layer_0[7706]; 
    assign out[536] = layer_0[3529] ^ layer_0[1595]; 
    assign out[537] = ~(layer_0[1770] ^ layer_0[1629]); 
    assign out[538] = layer_0[2161] ^ layer_0[6311]; 
    assign out[539] = ~layer_0[4407]; 
    assign out[540] = ~(layer_0[3889] ^ layer_0[468]); 
    assign out[541] = ~(layer_0[7976] ^ layer_0[5645]); 
    assign out[542] = layer_0[6026] ^ layer_0[2678]; 
    assign out[543] = layer_0[7634] & layer_0[3929]; 
    assign out[544] = ~layer_0[6107]; 
    assign out[545] = ~(layer_0[3522] ^ layer_0[6398]); 
    assign out[546] = layer_0[7239] & ~layer_0[2181]; 
    assign out[547] = layer_0[6644] ^ layer_0[542]; 
    assign out[548] = layer_0[4075] ^ layer_0[7535]; 
    assign out[549] = ~(layer_0[2010] ^ layer_0[2475]); 
    assign out[550] = layer_0[1117] & layer_0[7889]; 
    assign out[551] = layer_0[5568] ^ layer_0[4204]; 
    assign out[552] = ~(layer_0[5295] ^ layer_0[6972]); 
    assign out[553] = layer_0[7120]; 
    assign out[554] = layer_0[2919] ^ layer_0[12]; 
    assign out[555] = ~(layer_0[4316] ^ layer_0[7415]); 
    assign out[556] = layer_0[4415] ^ layer_0[4085]; 
    assign out[557] = layer_0[7522] & ~layer_0[2207]; 
    assign out[558] = layer_0[709] & ~layer_0[5659]; 
    assign out[559] = ~(layer_0[7082] ^ layer_0[1479]); 
    assign out[560] = ~(layer_0[2250] ^ layer_0[1775]); 
    assign out[561] = ~(layer_0[1797] & layer_0[6515]); 
    assign out[562] = ~layer_0[2200]; 
    assign out[563] = ~(layer_0[4473] ^ layer_0[653]); 
    assign out[564] = layer_0[2964] | layer_0[6301]; 
    assign out[565] = ~layer_0[3569]; 
    assign out[566] = ~(layer_0[7629] | layer_0[5475]); 
    assign out[567] = ~(layer_0[558] ^ layer_0[2929]); 
    assign out[568] = layer_0[4544]; 
    assign out[569] = layer_0[7426] ^ layer_0[4427]; 
    assign out[570] = ~(layer_0[2376] ^ layer_0[2154]); 
    assign out[571] = ~(layer_0[41] ^ layer_0[263]); 
    assign out[572] = layer_0[3114]; 
    assign out[573] = layer_0[5852] & ~layer_0[4680]; 
    assign out[574] = ~layer_0[7290]; 
    assign out[575] = layer_0[5221] | layer_0[6784]; 
    assign out[576] = layer_0[6004] | layer_0[4814]; 
    assign out[577] = layer_0[7815] ^ layer_0[6446]; 
    assign out[578] = layer_0[7900] ^ layer_0[1230]; 
    assign out[579] = ~(layer_0[5564] ^ layer_0[877]); 
    assign out[580] = layer_0[2685] & layer_0[2046]; 
    assign out[581] = ~layer_0[7179]; 
    assign out[582] = layer_0[222] ^ layer_0[1451]; 
    assign out[583] = layer_0[3431] ^ layer_0[899]; 
    assign out[584] = layer_0[6833] & ~layer_0[1094]; 
    assign out[585] = layer_0[7951] ^ layer_0[761]; 
    assign out[586] = layer_0[986] & ~layer_0[4854]; 
    assign out[587] = layer_0[4630] & ~layer_0[3931]; 
    assign out[588] = layer_0[2281] & ~layer_0[3717]; 
    assign out[589] = layer_0[5149]; 
    assign out[590] = ~(layer_0[815] & layer_0[377]); 
    assign out[591] = ~(layer_0[78] | layer_0[3001]); 
    assign out[592] = ~layer_0[4883]; 
    assign out[593] = layer_0[3837] & layer_0[5535]; 
    assign out[594] = layer_0[3947]; 
    assign out[595] = layer_0[5246] ^ layer_0[399]; 
    assign out[596] = layer_0[3539] | layer_0[7008]; 
    assign out[597] = layer_0[1197] ^ layer_0[6487]; 
    assign out[598] = ~(layer_0[7214] ^ layer_0[7950]); 
    assign out[599] = ~(layer_0[6355] ^ layer_0[705]); 
    assign out[600] = layer_0[4281]; 
    assign out[601] = ~layer_0[6258]; 
    assign out[602] = layer_0[5758] & ~layer_0[944]; 
    assign out[603] = layer_0[2517]; 
    assign out[604] = layer_0[7986] & ~layer_0[2372]; 
    assign out[605] = ~(layer_0[4869] ^ layer_0[328]); 
    assign out[606] = ~layer_0[5218]; 
    assign out[607] = layer_0[7399]; 
    assign out[608] = layer_0[1358] & layer_0[6312]; 
    assign out[609] = ~layer_0[651]; 
    assign out[610] = layer_0[1234] | layer_0[2662]; 
    assign out[611] = layer_0[4283] ^ layer_0[2218]; 
    assign out[612] = layer_0[4083] & ~layer_0[3401]; 
    assign out[613] = layer_0[206] ^ layer_0[1289]; 
    assign out[614] = ~layer_0[2319]; 
    assign out[615] = layer_0[7029] & layer_0[3356]; 
    assign out[616] = ~(layer_0[5410] | layer_0[4696]); 
    assign out[617] = ~layer_0[2814] | (layer_0[2814] & layer_0[6413]); 
    assign out[618] = ~(layer_0[3437] ^ layer_0[6361]); 
    assign out[619] = ~(layer_0[1065] ^ layer_0[5305]); 
    assign out[620] = ~layer_0[7278]; 
    assign out[621] = layer_0[5207] & layer_0[2398]; 
    assign out[622] = layer_0[4994]; 
    assign out[623] = ~(layer_0[42] ^ layer_0[5236]); 
    assign out[624] = layer_0[7031] ^ layer_0[3826]; 
    assign out[625] = ~(layer_0[7813] ^ layer_0[4383]); 
    assign out[626] = ~(layer_0[1170] ^ layer_0[1940]); 
    assign out[627] = layer_0[5283]; 
    assign out[628] = layer_0[6204] ^ layer_0[7943]; 
    assign out[629] = layer_0[5579] ^ layer_0[728]; 
    assign out[630] = ~(layer_0[744] | layer_0[4516]); 
    assign out[631] = ~(layer_0[7743] ^ layer_0[5794]); 
    assign out[632] = ~layer_0[4566]; 
    assign out[633] = layer_0[2641] | layer_0[4237]; 
    assign out[634] = layer_0[2644] ^ layer_0[2674]; 
    assign out[635] = ~(layer_0[4692] | layer_0[2396]); 
    assign out[636] = layer_0[74] ^ layer_0[5422]; 
    assign out[637] = ~layer_0[1474] | (layer_0[1474] & layer_0[1286]); 
    assign out[638] = layer_0[3896] ^ layer_0[3963]; 
    assign out[639] = ~(layer_0[7127] ^ layer_0[5279]); 
    assign out[640] = layer_0[6348]; 
    assign out[641] = layer_0[3520] ^ layer_0[5790]; 
    assign out[642] = layer_0[6866]; 
    assign out[643] = ~(layer_0[6245] ^ layer_0[3713]); 
    assign out[644] = layer_0[2232] & ~layer_0[2634]; 
    assign out[645] = ~(layer_0[1176] ^ layer_0[111]); 
    assign out[646] = layer_0[2351] ^ layer_0[5609]; 
    assign out[647] = layer_0[7389]; 
    assign out[648] = layer_0[1853]; 
    assign out[649] = layer_0[350] & ~layer_0[1863]; 
    assign out[650] = layer_0[7737]; 
    assign out[651] = layer_0[5552] & ~layer_0[3665]; 
    assign out[652] = ~(layer_0[4330] ^ layer_0[5292]); 
    assign out[653] = layer_0[2669]; 
    assign out[654] = layer_0[5101]; 
    assign out[655] = layer_0[2546] | layer_0[3351]; 
    assign out[656] = layer_0[1191]; 
    assign out[657] = ~(layer_0[4446] ^ layer_0[5700]); 
    assign out[658] = ~layer_0[1229] | (layer_0[6183] & layer_0[1229]); 
    assign out[659] = ~layer_0[1262]; 
    assign out[660] = layer_0[7532]; 
    assign out[661] = layer_0[298]; 
    assign out[662] = ~layer_0[7617] | (layer_0[6613] & layer_0[7617]); 
    assign out[663] = ~layer_0[1259] | (layer_0[1259] & layer_0[4658]); 
    assign out[664] = layer_0[2837] & ~layer_0[65]; 
    assign out[665] = ~(layer_0[836] ^ layer_0[3153]); 
    assign out[666] = ~layer_0[3902]; 
    assign out[667] = ~(layer_0[3373] ^ layer_0[4800]); 
    assign out[668] = layer_0[2113] | layer_0[5234]; 
    assign out[669] = ~(layer_0[2587] ^ layer_0[5359]); 
    assign out[670] = layer_0[2374] | layer_0[7061]; 
    assign out[671] = ~layer_0[6824]; 
    assign out[672] = layer_0[1604] ^ layer_0[604]; 
    assign out[673] = ~layer_0[7805]; 
    assign out[674] = ~(layer_0[1685] & layer_0[5146]); 
    assign out[675] = layer_0[2675]; 
    assign out[676] = ~(layer_0[3500] ^ layer_0[4708]); 
    assign out[677] = layer_0[2969] ^ layer_0[56]; 
    assign out[678] = layer_0[2679] ^ layer_0[6594]; 
    assign out[679] = ~layer_0[2681]; 
    assign out[680] = ~layer_0[5864]; 
    assign out[681] = layer_0[966] ^ layer_0[141]; 
    assign out[682] = layer_0[831] & layer_0[3734]; 
    assign out[683] = layer_0[1122] ^ layer_0[2846]; 
    assign out[684] = ~layer_0[7327] | (layer_0[952] & layer_0[7327]); 
    assign out[685] = layer_0[2744] ^ layer_0[7214]; 
    assign out[686] = ~layer_0[91]; 
    assign out[687] = layer_0[3676] | layer_0[6279]; 
    assign out[688] = ~layer_0[7134]; 
    assign out[689] = ~(layer_0[235] ^ layer_0[3867]); 
    assign out[690] = layer_0[5467]; 
    assign out[691] = ~layer_0[7557] | (layer_0[7557] & layer_0[2898]); 
    assign out[692] = ~layer_0[4397]; 
    assign out[693] = ~(layer_0[5867] ^ layer_0[5118]); 
    assign out[694] = layer_0[6565] ^ layer_0[5249]; 
    assign out[695] = layer_0[6053] & layer_0[7340]; 
    assign out[696] = ~layer_0[5882] | (layer_0[5882] & layer_0[7217]); 
    assign out[697] = ~(layer_0[2839] ^ layer_0[7208]); 
    assign out[698] = layer_0[886] | layer_0[5940]; 
    assign out[699] = ~layer_0[3418]; 
    assign out[700] = ~layer_0[5906] | (layer_0[5906] & layer_0[140]); 
    assign out[701] = layer_0[766] ^ layer_0[5484]; 
    assign out[702] = ~(layer_0[5747] ^ layer_0[1866]); 
    assign out[703] = ~(layer_0[3428] ^ layer_0[1937]); 
    assign out[704] = layer_0[3377] & ~layer_0[2667]; 
    assign out[705] = layer_0[4558] ^ layer_0[4259]; 
    assign out[706] = ~(layer_0[299] ^ layer_0[4637]); 
    assign out[707] = layer_0[7529] & ~layer_0[4138]; 
    assign out[708] = layer_0[2091] & ~layer_0[1610]; 
    assign out[709] = ~(layer_0[3937] ^ layer_0[3013]); 
    assign out[710] = layer_0[5222] ^ layer_0[872]; 
    assign out[711] = layer_0[4582] ^ layer_0[4735]; 
    assign out[712] = layer_0[13] | layer_0[589]; 
    assign out[713] = layer_0[5002] & ~layer_0[131]; 
    assign out[714] = layer_0[5486]; 
    assign out[715] = ~layer_0[1644] | (layer_0[5479] & layer_0[1644]); 
    assign out[716] = layer_0[3842] & layer_0[1276]; 
    assign out[717] = layer_0[2180] & ~layer_0[4478]; 
    assign out[718] = layer_0[797] ^ layer_0[333]; 
    assign out[719] = ~(layer_0[5873] ^ layer_0[39]); 
    assign out[720] = ~(layer_0[3794] ^ layer_0[4123]); 
    assign out[721] = layer_0[671] ^ layer_0[3012]; 
    assign out[722] = ~(layer_0[4258] ^ layer_0[1539]); 
    assign out[723] = layer_0[1315] & ~layer_0[5781]; 
    assign out[724] = layer_0[6379] & layer_0[4071]; 
    assign out[725] = layer_0[4733]; 
    assign out[726] = ~layer_0[1532]; 
    assign out[727] = ~(layer_0[5658] ^ layer_0[5611]); 
    assign out[728] = ~(layer_0[3922] ^ layer_0[652]); 
    assign out[729] = layer_0[1077]; 
    assign out[730] = layer_0[4239] ^ layer_0[7467]; 
    assign out[731] = layer_0[2130] & ~layer_0[2877]; 
    assign out[732] = layer_0[2876] & ~layer_0[7912]; 
    assign out[733] = ~(layer_0[5942] | layer_0[3802]); 
    assign out[734] = layer_0[4545] & ~layer_0[7996]; 
    assign out[735] = layer_0[7499]; 
    assign out[736] = ~(layer_0[2059] ^ layer_0[6505]); 
    assign out[737] = ~layer_0[5736] | (layer_0[4700] & layer_0[5736]); 
    assign out[738] = layer_0[4556]; 
    assign out[739] = layer_0[6584] & ~layer_0[4558]; 
    assign out[740] = ~(layer_0[7] ^ layer_0[4405]); 
    assign out[741] = ~(layer_0[4443] | layer_0[6930]); 
    assign out[742] = layer_0[6676] & ~layer_0[6136]; 
    assign out[743] = ~(layer_0[90] ^ layer_0[4154]); 
    assign out[744] = ~layer_0[6084] | (layer_0[40] & layer_0[6084]); 
    assign out[745] = ~layer_0[5127]; 
    assign out[746] = layer_0[6366] & ~layer_0[1883]; 
    assign out[747] = layer_0[4112] ^ layer_0[6045]; 
    assign out[748] = ~(layer_0[7304] ^ layer_0[5593]); 
    assign out[749] = ~(layer_0[5337] & layer_0[3789]); 
    assign out[750] = ~(layer_0[959] ^ layer_0[2492]); 
    assign out[751] = ~(layer_0[1649] ^ layer_0[5333]); 
    assign out[752] = layer_0[7434]; 
    assign out[753] = ~layer_0[6288]; 
    assign out[754] = layer_0[2808] ^ layer_0[2831]; 
    assign out[755] = layer_0[7476] ^ layer_0[240]; 
    assign out[756] = layer_0[702]; 
    assign out[757] = layer_0[7028] ^ layer_0[6334]; 
    assign out[758] = layer_0[5565] & ~layer_0[6047]; 
    assign out[759] = layer_0[7457]; 
    assign out[760] = layer_0[5194]; 
    assign out[761] = ~(layer_0[2322] ^ layer_0[3548]); 
    assign out[762] = ~layer_0[7062] | (layer_0[3860] & layer_0[7062]); 
    assign out[763] = ~(layer_0[5036] | layer_0[1001]); 
    assign out[764] = layer_0[7085]; 
    assign out[765] = ~(layer_0[429] ^ layer_0[5229]); 
    assign out[766] = layer_0[1232] ^ layer_0[1058]; 
    assign out[767] = layer_0[5293] & ~layer_0[3330]; 
    assign out[768] = layer_0[1068] ^ layer_0[1163]; 
    assign out[769] = ~(layer_0[1136] ^ layer_0[2637]); 
    assign out[770] = ~layer_0[4781]; 
    assign out[771] = layer_0[4329] ^ layer_0[2793]; 
    assign out[772] = layer_0[5685] ^ layer_0[7418]; 
    assign out[773] = ~(layer_0[763] ^ layer_0[5306]); 
    assign out[774] = layer_0[5301] ^ layer_0[3928]; 
    assign out[775] = layer_0[5121] ^ layer_0[2242]; 
    assign out[776] = layer_0[180] & ~layer_0[6925]; 
    assign out[777] = ~(layer_0[3723] ^ layer_0[3954]); 
    assign out[778] = ~layer_0[940]; 
    assign out[779] = ~(layer_0[1522] ^ layer_0[6865]); 
    assign out[780] = layer_0[1349] & layer_0[2478]; 
    assign out[781] = ~(layer_0[6822] ^ layer_0[3505]); 
    assign out[782] = layer_0[3004]; 
    assign out[783] = ~layer_0[4955] | (layer_0[1088] & layer_0[4955]); 
    assign out[784] = layer_0[4309] ^ layer_0[3687]; 
    assign out[785] = layer_0[99] & ~layer_0[5840]; 
    assign out[786] = layer_0[5709] ^ layer_0[4707]; 
    assign out[787] = ~layer_0[6778] | (layer_0[3560] & layer_0[6778]); 
    assign out[788] = layer_0[6583] ^ layer_0[4580]; 
    assign out[789] = layer_0[5415] | layer_0[4028]; 
    assign out[790] = ~(layer_0[6904] ^ layer_0[5077]); 
    assign out[791] = ~layer_0[4614]; 
    assign out[792] = layer_0[2220] & ~layer_0[1743]; 
    assign out[793] = 1'b1; 
    assign out[794] = ~layer_0[6948]; 
    assign out[795] = ~(layer_0[2427] ^ layer_0[1528]); 
    assign out[796] = layer_0[2937] ^ layer_0[6320]; 
    assign out[797] = layer_0[6438] & ~layer_0[1794]; 
    assign out[798] = layer_0[720] ^ layer_0[3074]; 
    assign out[799] = layer_0[1647] & ~layer_0[4010]; 
    assign out[800] = layer_0[7728] ^ layer_0[1870]; 
    assign out[801] = ~(layer_0[4528] ^ layer_0[2495]); 
    assign out[802] = ~(layer_0[1822] ^ layer_0[1885]); 
    assign out[803] = ~layer_0[3936]; 
    assign out[804] = layer_0[6908] & ~layer_0[200]; 
    assign out[805] = layer_0[5026] ^ layer_0[7551]; 
    assign out[806] = layer_0[4636]; 
    assign out[807] = layer_0[4959] & ~layer_0[6615]; 
    assign out[808] = layer_0[5981]; 
    assign out[809] = layer_0[3703] ^ layer_0[7074]; 
    assign out[810] = ~layer_0[3080]; 
    assign out[811] = layer_0[5436] ^ layer_0[7833]; 
    assign out[812] = ~(layer_0[5509] | layer_0[95]); 
    assign out[813] = ~layer_0[6668] | (layer_0[6668] & layer_0[929]); 
    assign out[814] = layer_0[1662]; 
    assign out[815] = ~layer_0[7075]; 
    assign out[816] = ~(layer_0[4191] ^ layer_0[1683]); 
    assign out[817] = layer_0[2763] ^ layer_0[6484]; 
    assign out[818] = layer_0[6414] & layer_0[6226]; 
    assign out[819] = ~layer_0[6945]; 
    assign out[820] = layer_0[1871] ^ layer_0[5834]; 
    assign out[821] = layer_0[6664] ^ layer_0[3946]; 
    assign out[822] = layer_0[2774]; 
    assign out[823] = layer_0[2389] | layer_0[6625]; 
    assign out[824] = ~(layer_0[1274] ^ layer_0[1772]); 
    assign out[825] = layer_0[225] & ~layer_0[2223]; 
    assign out[826] = layer_0[1654]; 
    assign out[827] = ~layer_0[2375]; 
    assign out[828] = layer_0[2043] ^ layer_0[1163]; 
    assign out[829] = ~layer_0[945] | (layer_0[945] & layer_0[155]); 
    assign out[830] = ~(layer_0[6185] ^ layer_0[166]); 
    assign out[831] = layer_0[7002] ^ layer_0[1625]; 
    assign out[832] = ~layer_0[3623]; 
    assign out[833] = layer_0[6228]; 
    assign out[834] = ~(layer_0[1265] & layer_0[6]); 
    assign out[835] = layer_0[3247] ^ layer_0[1461]; 
    assign out[836] = layer_0[5544] ^ layer_0[5517]; 
    assign out[837] = layer_0[2548]; 
    assign out[838] = layer_0[2963]; 
    assign out[839] = ~layer_0[2970]; 
    assign out[840] = ~layer_0[5063]; 
    assign out[841] = ~layer_0[3494]; 
    assign out[842] = ~(layer_0[2664] | layer_0[6574]); 
    assign out[843] = ~layer_0[5431] | (layer_0[4783] & layer_0[5431]); 
    assign out[844] = layer_0[2725] | layer_0[150]; 
    assign out[845] = ~layer_0[133]; 
    assign out[846] = layer_0[5358] ^ layer_0[4374]; 
    assign out[847] = ~(layer_0[5763] ^ layer_0[3606]); 
    assign out[848] = layer_0[6226]; 
    assign out[849] = ~layer_0[292]; 
    assign out[850] = layer_0[5408] ^ layer_0[3499]; 
    assign out[851] = ~(layer_0[2419] ^ layer_0[2575]); 
    assign out[852] = layer_0[320] ^ layer_0[2403]; 
    assign out[853] = ~layer_0[3127]; 
    assign out[854] = layer_0[3918]; 
    assign out[855] = ~(layer_0[6704] ^ layer_0[6090]); 
    assign out[856] = ~(layer_0[5217] & layer_0[5435]); 
    assign out[857] = ~(layer_0[5549] ^ layer_0[4786]); 
    assign out[858] = layer_0[1800] ^ layer_0[2827]; 
    assign out[859] = ~layer_0[1445]; 
    assign out[860] = ~(layer_0[3390] ^ layer_0[7832]); 
    assign out[861] = layer_0[3073] ^ layer_0[974]; 
    assign out[862] = layer_0[4507] & ~layer_0[960]; 
    assign out[863] = layer_0[4507]; 
    assign out[864] = ~(layer_0[4940] ^ layer_0[4344]); 
    assign out[865] = layer_0[2239] & ~layer_0[717]; 
    assign out[866] = ~(layer_0[7796] ^ layer_0[555]); 
    assign out[867] = layer_0[3921] & ~layer_0[2667]; 
    assign out[868] = ~(layer_0[1586] ^ layer_0[3878]); 
    assign out[869] = ~(layer_0[7060] ^ layer_0[7636]); 
    assign out[870] = layer_0[3140] & layer_0[2739]; 
    assign out[871] = ~layer_0[5860]; 
    assign out[872] = layer_0[2830] ^ layer_0[7007]; 
    assign out[873] = ~(layer_0[3617] ^ layer_0[7190]); 
    assign out[874] = ~(layer_0[3398] & layer_0[1004]); 
    assign out[875] = layer_0[6797] ^ layer_0[5660]; 
    assign out[876] = ~(layer_0[4321] ^ layer_0[5808]); 
    assign out[877] = layer_0[5758]; 
    assign out[878] = layer_0[6945]; 
    assign out[879] = layer_0[1512] ^ layer_0[656]; 
    assign out[880] = layer_0[882] ^ layer_0[822]; 
    assign out[881] = layer_0[5908] ^ layer_0[1786]; 
    assign out[882] = layer_0[5625] ^ layer_0[1401]; 
    assign out[883] = ~(layer_0[4963] ^ layer_0[4957]); 
    assign out[884] = layer_0[7666] | layer_0[7162]; 
    assign out[885] = layer_0[6597] ^ layer_0[3254]; 
    assign out[886] = ~(layer_0[1160] | layer_0[4912]); 
    assign out[887] = layer_0[3568] | layer_0[5882]; 
    assign out[888] = layer_0[2422] ^ layer_0[1534]; 
    assign out[889] = layer_0[5154] & layer_0[854]; 
    assign out[890] = ~(layer_0[2220] & layer_0[2654]); 
    assign out[891] = ~layer_0[1035] | (layer_0[2302] & layer_0[1035]); 
    assign out[892] = ~layer_0[6684]; 
    assign out[893] = layer_0[4030]; 
    assign out[894] = layer_0[1630]; 
    assign out[895] = layer_0[2772] | layer_0[7408]; 
    assign out[896] = layer_0[917] & layer_0[869]; 
    assign out[897] = ~(layer_0[7273] ^ layer_0[3134]); 
    assign out[898] = layer_0[3456] & ~layer_0[6286]; 
    assign out[899] = ~(layer_0[4018] | layer_0[7615]); 
    assign out[900] = layer_0[2815] ^ layer_0[5191]; 
    assign out[901] = layer_0[1962] ^ layer_0[6524]; 
    assign out[902] = layer_0[6871] ^ layer_0[4340]; 
    assign out[903] = ~layer_0[1908]; 
    assign out[904] = ~layer_0[4689]; 
    assign out[905] = ~(layer_0[5741] ^ layer_0[1460]); 
    assign out[906] = layer_0[4706] & layer_0[2418]; 
    assign out[907] = layer_0[1132]; 
    assign out[908] = layer_0[6006] ^ layer_0[355]; 
    assign out[909] = layer_0[6058] ^ layer_0[2735]; 
    assign out[910] = layer_0[697] ^ layer_0[5639]; 
    assign out[911] = layer_0[6748] & ~layer_0[6581]; 
    assign out[912] = ~layer_0[7432]; 
    assign out[913] = layer_0[1579] ^ layer_0[3489]; 
    assign out[914] = layer_0[773] ^ layer_0[6278]; 
    assign out[915] = layer_0[4257]; 
    assign out[916] = layer_0[6170]; 
    assign out[917] = ~layer_0[5883] | (layer_0[5883] & layer_0[5971]); 
    assign out[918] = layer_0[861] & layer_0[3093]; 
    assign out[919] = layer_0[274] & layer_0[4080]; 
    assign out[920] = layer_0[3751] & layer_0[1679]; 
    assign out[921] = ~(layer_0[3392] ^ layer_0[5526]); 
    assign out[922] = ~(layer_0[2205] ^ layer_0[129]); 
    assign out[923] = ~layer_0[6423]; 
    assign out[924] = ~(layer_0[7337] & layer_0[1211]); 
    assign out[925] = layer_0[2574] & layer_0[6193]; 
    assign out[926] = layer_0[152]; 
    assign out[927] = ~(layer_0[3993] & layer_0[2900]); 
    assign out[928] = layer_0[7774] ^ layer_0[1608]; 
    assign out[929] = layer_0[2571]; 
    assign out[930] = layer_0[4697]; 
    assign out[931] = layer_0[7732] ^ layer_0[5816]; 
    assign out[932] = layer_0[5115] ^ layer_0[7435]; 
    assign out[933] = layer_0[3035] ^ layer_0[7921]; 
    assign out[934] = layer_0[5844] ^ layer_0[2482]; 
    assign out[935] = layer_0[4114] ^ layer_0[1227]; 
    assign out[936] = layer_0[2683] & ~layer_0[2665]; 
    assign out[937] = layer_0[3747] ^ layer_0[6598]; 
    assign out[938] = ~layer_0[4410]; 
    assign out[939] = ~layer_0[2292] | (layer_0[2292] & layer_0[3110]); 
    assign out[940] = layer_0[620] & ~layer_0[2190]; 
    assign out[941] = layer_0[5623] & layer_0[1298]; 
    assign out[942] = ~(layer_0[4617] | layer_0[5178]); 
    assign out[943] = layer_0[5868] ^ layer_0[5421]; 
    assign out[944] = layer_0[7713] & ~layer_0[7795]; 
    assign out[945] = ~(layer_0[3996] ^ layer_0[4137]); 
    assign out[946] = layer_0[5069] ^ layer_0[4542]; 
    assign out[947] = layer_0[2328] & ~layer_0[278]; 
    assign out[948] = layer_0[7572]; 
    assign out[949] = layer_0[1036] & layer_0[2962]; 
    assign out[950] = layer_0[6725]; 
    assign out[951] = layer_0[5887] ^ layer_0[4672]; 
    assign out[952] = ~(layer_0[2817] ^ layer_0[1339]); 
    assign out[953] = layer_0[7307] & ~layer_0[2318]; 
    assign out[954] = layer_0[2784]; 
    assign out[955] = layer_0[7844]; 
    assign out[956] = layer_0[7106] & ~layer_0[6545]; 
    assign out[957] = layer_0[7747] ^ layer_0[4698]; 
    assign out[958] = layer_0[4337] | layer_0[4251]; 
    assign out[959] = layer_0[1672] ^ layer_0[4800]; 
    assign out[960] = ~layer_0[6717] | (layer_0[2645] & layer_0[6717]); 
    assign out[961] = layer_0[7594] & layer_0[3668]; 
    assign out[962] = layer_0[6150] & ~layer_0[5606]; 
    assign out[963] = ~layer_0[677]; 
    assign out[964] = ~(layer_0[3659] | layer_0[4136]); 
    assign out[965] = layer_0[7407] & ~layer_0[621]; 
    assign out[966] = layer_0[5580] & ~layer_0[1696]; 
    assign out[967] = layer_0[5154] & layer_0[2493]; 
    assign out[968] = ~(layer_0[496] ^ layer_0[895]); 
    assign out[969] = layer_0[1158] ^ layer_0[3958]; 
    assign out[970] = ~(layer_0[2992] ^ layer_0[659]); 
    assign out[971] = ~(layer_0[7145] ^ layer_0[1222]); 
    assign out[972] = layer_0[5848] ^ layer_0[3514]; 
    assign out[973] = layer_0[4228]; 
    assign out[974] = layer_0[3288] & ~layer_0[7395]; 
    assign out[975] = layer_0[7273]; 
    assign out[976] = ~layer_0[251]; 
    assign out[977] = layer_0[6529]; 
    assign out[978] = layer_0[3760] ^ layer_0[1352]; 
    assign out[979] = ~(layer_0[1977] ^ layer_0[5078]); 
    assign out[980] = layer_0[6982] ^ layer_0[3436]; 
    assign out[981] = ~(layer_0[1514] ^ layer_0[4667]); 
    assign out[982] = ~layer_0[2096]; 
    assign out[983] = ~(layer_0[5736] | layer_0[2709]); 
    assign out[984] = layer_0[7794] ^ layer_0[2588]; 
    assign out[985] = ~layer_0[296]; 
    assign out[986] = layer_0[6323]; 
    assign out[987] = ~(layer_0[4649] ^ layer_0[3192]); 
    assign out[988] = ~layer_0[6939]; 
    assign out[989] = layer_0[5116] ^ layer_0[1416]; 
    assign out[990] = layer_0[3391] ^ layer_0[1887]; 
    assign out[991] = layer_0[6575] ^ layer_0[2622]; 
    assign out[992] = ~(layer_0[2655] ^ layer_0[3990]); 
    assign out[993] = ~layer_0[3832]; 
    assign out[994] = ~(layer_0[427] ^ layer_0[4110]); 
    assign out[995] = ~(layer_0[3253] & layer_0[2381]); 
    assign out[996] = ~(layer_0[7978] & layer_0[3137]); 
    assign out[997] = ~layer_0[2818] | (layer_0[2818] & layer_0[2016]); 
    assign out[998] = ~layer_0[842]; 
    assign out[999] = layer_0[5646] ^ layer_0[938]; 
    assign out[1000] = ~layer_0[4629]; 
    assign out[1001] = ~layer_0[2602]; 
    assign out[1002] = layer_0[5345] ^ layer_0[6490]; 
    assign out[1003] = ~layer_0[582]; 
    assign out[1004] = ~(layer_0[6510] ^ layer_0[2222]); 
    assign out[1005] = ~layer_0[4251]; 
    assign out[1006] = ~(layer_0[7725] | layer_0[117]); 
    assign out[1007] = ~(layer_0[5062] ^ layer_0[4961]); 
    assign out[1008] = layer_0[2490] ^ layer_0[2843]; 
    assign out[1009] = ~layer_0[6663]; 
    assign out[1010] = ~layer_0[7441]; 
    assign out[1011] = ~layer_0[2303]; 
    assign out[1012] = ~layer_0[3041]; 
    assign out[1013] = ~(layer_0[4426] ^ layer_0[289]); 
    assign out[1014] = layer_0[5890] ^ layer_0[2825]; 
    assign out[1015] = ~(layer_0[3846] ^ layer_0[3800]); 
    assign out[1016] = layer_0[5214] & layer_0[6242]; 
    assign out[1017] = layer_0[3555]; 
    assign out[1018] = ~(layer_0[5878] ^ layer_0[5753]); 
    assign out[1019] = ~(layer_0[4522] ^ layer_0[7033]); 
    assign out[1020] = layer_0[4108] & layer_0[1306]; 
    assign out[1021] = ~layer_0[1730]; 
    assign out[1022] = layer_0[5654] ^ layer_0[5853]; 
    assign out[1023] = layer_0[5283] ^ layer_0[7813]; 
    assign out[1024] = layer_0[1801] ^ layer_0[1391]; 
    assign out[1025] = layer_0[2236] | layer_0[4087]; 
    assign out[1026] = ~(layer_0[7245] ^ layer_0[5766]); 
    assign out[1027] = layer_0[3696] ^ layer_0[7767]; 
    assign out[1028] = ~layer_0[6626]; 
    assign out[1029] = layer_0[5600] ^ layer_0[4260]; 
    assign out[1030] = ~(layer_0[7072] ^ layer_0[5533]); 
    assign out[1031] = ~layer_0[7025]; 
    assign out[1032] = layer_0[1485] ^ layer_0[4651]; 
    assign out[1033] = layer_0[5123] ^ layer_0[579]; 
    assign out[1034] = layer_0[4664] ^ layer_0[6661]; 
    assign out[1035] = layer_0[7895] & ~layer_0[4815]; 
    assign out[1036] = layer_0[7688] ^ layer_0[5237]; 
    assign out[1037] = ~(layer_0[730] | layer_0[1319]); 
    assign out[1038] = layer_0[7158] ^ layer_0[5353]; 
    assign out[1039] = layer_0[7437] ^ layer_0[550]; 
    assign out[1040] = layer_0[5324] ^ layer_0[4489]; 
    assign out[1041] = ~layer_0[1092]; 
    assign out[1042] = ~layer_0[1347] | (layer_0[344] & layer_0[1347]); 
    assign out[1043] = ~layer_0[1562] | (layer_0[2529] & layer_0[1562]); 
    assign out[1044] = layer_0[1948]; 
    assign out[1045] = layer_0[7421] & ~layer_0[4166]; 
    assign out[1046] = layer_0[3956] ^ layer_0[4298]; 
    assign out[1047] = layer_0[4987]; 
    assign out[1048] = ~layer_0[5049] | (layer_0[5049] & layer_0[2057]); 
    assign out[1049] = ~(layer_0[5145] ^ layer_0[3838]); 
    assign out[1050] = layer_0[6567]; 
    assign out[1051] = ~(layer_0[2585] ^ layer_0[4428]); 
    assign out[1052] = ~(layer_0[2979] ^ layer_0[619]); 
    assign out[1053] = layer_0[6307] ^ layer_0[2359]; 
    assign out[1054] = ~layer_0[1909]; 
    assign out[1055] = ~(layer_0[115] | layer_0[5227]); 
    assign out[1056] = layer_0[218]; 
    assign out[1057] = ~layer_0[517]; 
    assign out[1058] = layer_0[6122]; 
    assign out[1059] = layer_0[4765] & ~layer_0[6472]; 
    assign out[1060] = layer_0[7320] ^ layer_0[2921]; 
    assign out[1061] = ~(layer_0[7989] ^ layer_0[1728]); 
    assign out[1062] = layer_0[5618] | layer_0[1584]; 
    assign out[1063] = layer_0[120]; 
    assign out[1064] = ~layer_0[4220] | (layer_0[4220] & layer_0[2016]); 
    assign out[1065] = ~layer_0[216]; 
    assign out[1066] = layer_0[2155] ^ layer_0[3362]; 
    assign out[1067] = layer_0[6254] ^ layer_0[7378]; 
    assign out[1068] = layer_0[7521] ^ layer_0[1873]; 
    assign out[1069] = layer_0[533] ^ layer_0[5212]; 
    assign out[1070] = ~(layer_0[4447] ^ layer_0[1370]); 
    assign out[1071] = layer_0[3108] & ~layer_0[6320]; 
    assign out[1072] = layer_0[6111]; 
    assign out[1073] = ~(layer_0[2722] ^ layer_0[7948]); 
    assign out[1074] = layer_0[6758] ^ layer_0[6800]; 
    assign out[1075] = ~(layer_0[6580] ^ layer_0[7403]); 
    assign out[1076] = ~(layer_0[858] | layer_0[1916]); 
    assign out[1077] = ~layer_0[1664] | (layer_0[1664] & layer_0[7168]); 
    assign out[1078] = layer_0[1261]; 
    assign out[1079] = ~layer_0[4009] | (layer_0[4009] & layer_0[1415]); 
    assign out[1080] = ~(layer_0[615] & layer_0[2798]); 
    assign out[1081] = ~(layer_0[366] ^ layer_0[7616]); 
    assign out[1082] = layer_0[4767] & layer_0[4324]; 
    assign out[1083] = layer_0[313] ^ layer_0[4638]; 
    assign out[1084] = layer_0[723] ^ layer_0[7764]; 
    assign out[1085] = ~layer_0[4482]; 
    assign out[1086] = layer_0[4463]; 
    assign out[1087] = layer_0[7673] ^ layer_0[4444]; 
    assign out[1088] = layer_0[5507] ^ layer_0[7564]; 
    assign out[1089] = ~layer_0[7938]; 
    assign out[1090] = layer_0[2693] & layer_0[3091]; 
    assign out[1091] = layer_0[1101] ^ layer_0[2619]; 
    assign out[1092] = layer_0[7341] ^ layer_0[7217]; 
    assign out[1093] = layer_0[6546]; 
    assign out[1094] = layer_0[2341] ^ layer_0[7222]; 
    assign out[1095] = layer_0[3315] ^ layer_0[4917]; 
    assign out[1096] = ~(layer_0[4096] ^ layer_0[4593]); 
    assign out[1097] = layer_0[1677] & ~layer_0[4981]; 
    assign out[1098] = layer_0[2702] & layer_0[3518]; 
    assign out[1099] = ~(layer_0[2417] ^ layer_0[5164]); 
    assign out[1100] = ~layer_0[6831] | (layer_0[6831] & layer_0[5983]); 
    assign out[1101] = layer_0[2443] ^ layer_0[516]; 
    assign out[1102] = ~(layer_0[1137] ^ layer_0[1127]); 
    assign out[1103] = ~(layer_0[6315] & layer_0[1488]); 
    assign out[1104] = ~(layer_0[1212] ^ layer_0[6624]); 
    assign out[1105] = layer_0[6279] | layer_0[6556]; 
    assign out[1106] = layer_0[651] ^ layer_0[6460]; 
    assign out[1107] = ~(layer_0[786] ^ layer_0[5314]); 
    assign out[1108] = layer_0[7092] ^ layer_0[7576]; 
    assign out[1109] = ~(layer_0[2875] ^ layer_0[2450]); 
    assign out[1110] = ~(layer_0[1313] ^ layer_0[5340]); 
    assign out[1111] = ~layer_0[1044]; 
    assign out[1112] = ~(layer_0[1931] ^ layer_0[4249]); 
    assign out[1113] = layer_0[5411] ^ layer_0[684]; 
    assign out[1114] = layer_0[7372] ^ layer_0[2147]; 
    assign out[1115] = ~(layer_0[5208] ^ layer_0[3062]); 
    assign out[1116] = ~(layer_0[3998] & layer_0[6630]); 
    assign out[1117] = layer_0[7078] | layer_0[477]; 
    assign out[1118] = ~layer_0[1515] | (layer_0[1515] & layer_0[4299]); 
    assign out[1119] = layer_0[7603]; 
    assign out[1120] = ~(layer_0[5195] ^ layer_0[156]); 
    assign out[1121] = layer_0[1372] ^ layer_0[760]; 
    assign out[1122] = ~layer_0[1441]; 
    assign out[1123] = ~layer_0[3741] | (layer_0[1145] & layer_0[3741]); 
    assign out[1124] = layer_0[6003] ^ layer_0[802]; 
    assign out[1125] = layer_0[4856] ^ layer_0[2796]; 
    assign out[1126] = layer_0[3810] ^ layer_0[1047]; 
    assign out[1127] = ~(layer_0[5043] ^ layer_0[2736]); 
    assign out[1128] = ~(layer_0[7009] ^ layer_0[1380]); 
    assign out[1129] = ~(layer_0[2781] ^ layer_0[105]); 
    assign out[1130] = layer_0[3927] & layer_0[4763]; 
    assign out[1131] = ~(layer_0[7138] ^ layer_0[1718]); 
    assign out[1132] = ~(layer_0[4133] ^ layer_0[5216]); 
    assign out[1133] = ~(layer_0[2533] ^ layer_0[1527]); 
    assign out[1134] = layer_0[5472] ^ layer_0[3151]; 
    assign out[1135] = layer_0[3985] & ~layer_0[6801]; 
    assign out[1136] = layer_0[6761] ^ layer_0[7586]; 
    assign out[1137] = layer_0[5745] ^ layer_0[5955]; 
    assign out[1138] = layer_0[6934]; 
    assign out[1139] = ~layer_0[1355]; 
    assign out[1140] = ~layer_0[2785] | (layer_0[2785] & layer_0[6739]); 
    assign out[1141] = layer_0[3897] ^ layer_0[7578]; 
    assign out[1142] = layer_0[4818]; 
    assign out[1143] = layer_0[1029] ^ layer_0[3628]; 
    assign out[1144] = ~(layer_0[3782] ^ layer_0[6430]); 
    assign out[1145] = ~layer_0[5065]; 
    assign out[1146] = layer_0[4078] & layer_0[5097]; 
    assign out[1147] = layer_0[1055] & ~layer_0[4783]; 
    assign out[1148] = ~layer_0[1013]; 
    assign out[1149] = layer_0[4775] ^ layer_0[1179]; 
    assign out[1150] = layer_0[721] | layer_0[3335]; 
    assign out[1151] = layer_0[7457] ^ layer_0[1233]; 
    assign out[1152] = layer_0[7044] & ~layer_0[4362]; 
    assign out[1153] = layer_0[1657] ^ layer_0[4324]; 
    assign out[1154] = layer_0[2124] & ~layer_0[660]; 
    assign out[1155] = layer_0[5146] | layer_0[832]; 
    assign out[1156] = ~(layer_0[4684] ^ layer_0[1500]); 
    assign out[1157] = ~(layer_0[4641] ^ layer_0[4207]); 
    assign out[1158] = layer_0[2258] ^ layer_0[4983]; 
    assign out[1159] = layer_0[2731] ^ layer_0[186]; 
    assign out[1160] = ~(layer_0[3819] ^ layer_0[2710]); 
    assign out[1161] = layer_0[6958] | layer_0[746]; 
    assign out[1162] = ~(layer_0[5371] ^ layer_0[514]); 
    assign out[1163] = layer_0[283] & ~layer_0[4931]; 
    assign out[1164] = ~layer_0[3079]; 
    assign out[1165] = ~(layer_0[1308] | layer_0[6678]); 
    assign out[1166] = ~(layer_0[3839] ^ layer_0[4945]); 
    assign out[1167] = ~layer_0[5343] | (layer_0[5273] & layer_0[5343]); 
    assign out[1168] = layer_0[4307] ^ layer_0[3750]; 
    assign out[1169] = layer_0[3365] ^ layer_0[4772]; 
    assign out[1170] = ~(layer_0[7769] ^ layer_0[6218]); 
    assign out[1171] = ~layer_0[6316]; 
    assign out[1172] = layer_0[4741] | layer_0[767]; 
    assign out[1173] = layer_0[326] & ~layer_0[637]; 
    assign out[1174] = layer_0[2076] & layer_0[498]; 
    assign out[1175] = layer_0[4082] ^ layer_0[3694]; 
    assign out[1176] = ~(layer_0[7184] | layer_0[641]); 
    assign out[1177] = ~(layer_0[7546] ^ layer_0[5948]); 
    assign out[1178] = layer_0[4560] ^ layer_0[5727]; 
    assign out[1179] = ~(layer_0[5617] ^ layer_0[447]); 
    assign out[1180] = layer_0[5941] & ~layer_0[7042]; 
    assign out[1181] = ~layer_0[4858] | (layer_0[4858] & layer_0[908]); 
    assign out[1182] = ~layer_0[418]; 
    assign out[1183] = layer_0[5170] & ~layer_0[4718]; 
    assign out[1184] = layer_0[1384] ^ layer_0[5929]; 
    assign out[1185] = layer_0[6405] & ~layer_0[5560]; 
    assign out[1186] = layer_0[1701] & ~layer_0[4740]; 
    assign out[1187] = layer_0[2442] ^ layer_0[1130]; 
    assign out[1188] = ~(layer_0[7533] ^ layer_0[78]); 
    assign out[1189] = ~layer_0[1181]; 
    assign out[1190] = ~layer_0[4173] | (layer_0[7875] & layer_0[4173]); 
    assign out[1191] = ~layer_0[7427]; 
    assign out[1192] = ~(layer_0[1789] ^ layer_0[3648]); 
    assign out[1193] = layer_0[7516]; 
    assign out[1194] = ~(layer_0[4789] ^ layer_0[4556]); 
    assign out[1195] = ~layer_0[3297] | (layer_0[11] & layer_0[3297]); 
    assign out[1196] = layer_0[4913] ^ layer_0[38]; 
    assign out[1197] = layer_0[59] ^ layer_0[388]; 
    assign out[1198] = ~(layer_0[6070] & layer_0[5124]); 
    assign out[1199] = layer_0[2703]; 
    assign out[1200] = ~layer_0[3781]; 
    assign out[1201] = layer_0[724]; 
    assign out[1202] = layer_0[4477]; 
    assign out[1203] = ~(layer_0[6694] ^ layer_0[4380]); 
    assign out[1204] = ~(layer_0[5832] | layer_0[3633]); 
    assign out[1205] = ~(layer_0[3025] ^ layer_0[3142]); 
    assign out[1206] = ~(layer_0[4375] | layer_0[5940]); 
    assign out[1207] = ~(layer_0[102] ^ layer_0[5266]); 
    assign out[1208] = layer_0[3698] ^ layer_0[951]; 
    assign out[1209] = ~(layer_0[7592] ^ layer_0[1267]); 
    assign out[1210] = layer_0[6957] ^ layer_0[4820]; 
    assign out[1211] = ~(layer_0[3888] & layer_0[3526]); 
    assign out[1212] = ~(layer_0[4683] ^ layer_0[2488]); 
    assign out[1213] = layer_0[7421] ^ layer_0[3973]; 
    assign out[1214] = ~(layer_0[4819] ^ layer_0[7444]); 
    assign out[1215] = layer_0[6517]; 
    assign out[1216] = layer_0[3132] ^ layer_0[7005]; 
    assign out[1217] = ~(layer_0[6793] ^ layer_0[5406]); 
    assign out[1218] = ~(layer_0[2769] & layer_0[3515]); 
    assign out[1219] = ~layer_0[22] | (layer_0[22] & layer_0[7846]); 
    assign out[1220] = ~layer_0[3540]; 
    assign out[1221] = layer_0[5699] ^ layer_0[7280]; 
    assign out[1222] = ~(layer_0[6083] ^ layer_0[1461]); 
    assign out[1223] = layer_0[570] & ~layer_0[3435]; 
    assign out[1224] = ~(layer_0[7362] ^ layer_0[3202]); 
    assign out[1225] = ~(layer_0[7715] ^ layer_0[1067]); 
    assign out[1226] = layer_0[5365] ^ layer_0[6752]; 
    assign out[1227] = ~layer_0[4791]; 
    assign out[1228] = layer_0[2986] ^ layer_0[1072]; 
    assign out[1229] = layer_0[7174] & layer_0[6508]; 
    assign out[1230] = layer_0[3705] | layer_0[3113]; 
    assign out[1231] = ~(layer_0[3813] ^ layer_0[1991]); 
    assign out[1232] = layer_0[3879] & layer_0[3525]; 
    assign out[1233] = layer_0[3333] ^ layer_0[1310]; 
    assign out[1234] = layer_0[5910] | layer_0[5030]; 
    assign out[1235] = layer_0[6973] ^ layer_0[5323]; 
    assign out[1236] = layer_0[561] & layer_0[1305]; 
    assign out[1237] = ~(layer_0[4654] ^ layer_0[1952]); 
    assign out[1238] = ~layer_0[2180] | (layer_0[6416] & layer_0[2180]); 
    assign out[1239] = layer_0[319] | layer_0[5633]; 
    assign out[1240] = ~(layer_0[5425] | layer_0[2230]); 
    assign out[1241] = ~layer_0[2653]; 
    assign out[1242] = layer_0[3692] & ~layer_0[3870]; 
    assign out[1243] = ~layer_0[962]; 
    assign out[1244] = ~(layer_0[7748] ^ layer_0[2113]); 
    assign out[1245] = ~(layer_0[4946] ^ layer_0[2934]); 
    assign out[1246] = ~(layer_0[5400] ^ layer_0[3441]); 
    assign out[1247] = layer_0[6115]; 
    assign out[1248] = ~(layer_0[5742] | layer_0[3459]); 
    assign out[1249] = layer_0[1133]; 
    assign out[1250] = ~(layer_0[7560] | layer_0[5029]); 
    assign out[1251] = layer_0[3416] ^ layer_0[6836]; 
    assign out[1252] = layer_0[3977] ^ layer_0[6186]; 
    assign out[1253] = layer_0[7120] ^ layer_0[3778]; 
    assign out[1254] = ~layer_0[5449] | (layer_0[5449] & layer_0[6326]); 
    assign out[1255] = ~layer_0[7627] | (layer_0[3481] & layer_0[7627]); 
    assign out[1256] = layer_0[6703] ^ layer_0[5838]; 
    assign out[1257] = ~(layer_0[3057] & layer_0[7556]); 
    assign out[1258] = ~(layer_0[6133] ^ layer_0[2349]); 
    assign out[1259] = layer_0[1427] ^ layer_0[1755]; 
    assign out[1260] = layer_0[600] ^ layer_0[403]; 
    assign out[1261] = ~(layer_0[1676] ^ layer_0[2669]); 
    assign out[1262] = layer_0[4669] & layer_0[163]; 
    assign out[1263] = ~(layer_0[7158] ^ layer_0[4300]); 
    assign out[1264] = layer_0[3480] | layer_0[4703]; 
    assign out[1265] = ~(layer_0[6453] ^ layer_0[1437]); 
    assign out[1266] = layer_0[7891] ^ layer_0[5897]; 
    assign out[1267] = layer_0[904]; 
    assign out[1268] = ~(layer_0[7567] ^ layer_0[5259]); 
    assign out[1269] = ~(layer_0[6821] & layer_0[890]); 
    assign out[1270] = layer_0[6814] & layer_0[6718]; 
    assign out[1271] = ~(layer_0[4925] ^ layer_0[3875]); 
    assign out[1272] = layer_0[2883] ^ layer_0[5691]; 
    assign out[1273] = ~(layer_0[6737] | layer_0[1104]); 
    assign out[1274] = layer_0[1264] ^ layer_0[3755]; 
    assign out[1275] = layer_0[4590] ^ layer_0[4625]; 
    assign out[1276] = ~(layer_0[3358] ^ layer_0[7860]); 
    assign out[1277] = ~(layer_0[2233] | layer_0[6631]); 
    assign out[1278] = ~layer_0[7071] | (layer_0[3636] & layer_0[7071]); 
    assign out[1279] = layer_0[6587]; 
    assign out[1280] = layer_0[7168] & ~layer_0[2993]; 
    assign out[1281] = ~(layer_0[3380] ^ layer_0[5308]); 
    assign out[1282] = layer_0[2305] & ~layer_0[7007]; 
    assign out[1283] = ~layer_0[3961]; 
    assign out[1284] = layer_0[866] & ~layer_0[3296]; 
    assign out[1285] = layer_0[1447] & ~layer_0[5963]; 
    assign out[1286] = layer_0[4730] ^ layer_0[437]; 
    assign out[1287] = ~layer_0[4341]; 
    assign out[1288] = ~(layer_0[996] ^ layer_0[5411]); 
    assign out[1289] = ~(layer_0[1838] ^ layer_0[1702]); 
    assign out[1290] = ~layer_0[1250]; 
    assign out[1291] = layer_0[6051] ^ layer_0[3573]; 
    assign out[1292] = ~(layer_0[2397] ^ layer_0[4220]); 
    assign out[1293] = layer_0[4525] & ~layer_0[5295]; 
    assign out[1294] = layer_0[3430] ^ layer_0[6638]; 
    assign out[1295] = layer_0[4523]; 
    assign out[1296] = layer_0[1162] ^ layer_0[1745]; 
    assign out[1297] = layer_0[564] ^ layer_0[5275]; 
    assign out[1298] = ~(layer_0[3893] ^ layer_0[3970]); 
    assign out[1299] = layer_0[422] ^ layer_0[2423]; 
    assign out[1300] = layer_0[1684] ^ layer_0[2445]; 
    assign out[1301] = ~layer_0[6621] | (layer_0[6621] & layer_0[6496]); 
    assign out[1302] = layer_0[2489] ^ layer_0[6134]; 
    assign out[1303] = layer_0[5506] ^ layer_0[7653]; 
    assign out[1304] = layer_0[3167] ^ layer_0[1992]; 
    assign out[1305] = ~(layer_0[915] ^ layer_0[2138]); 
    assign out[1306] = ~(layer_0[3015] | layer_0[686]); 
    assign out[1307] = ~(layer_0[3324] ^ layer_0[2933]); 
    assign out[1308] = ~(layer_0[4027] ^ layer_0[887]); 
    assign out[1309] = layer_0[2980] ^ layer_0[302]; 
    assign out[1310] = layer_0[3223] ^ layer_0[3627]; 
    assign out[1311] = layer_0[7170] ^ layer_0[5117]; 
    assign out[1312] = layer_0[5450] ^ layer_0[583]; 
    assign out[1313] = ~(layer_0[2945] ^ layer_0[5462]); 
    assign out[1314] = ~(layer_0[2032] ^ layer_0[3191]); 
    assign out[1315] = ~(layer_0[856] & layer_0[4095]); 
    assign out[1316] = ~layer_0[2650]; 
    assign out[1317] = ~(layer_0[5182] ^ layer_0[3943]); 
    assign out[1318] = ~(layer_0[6922] ^ layer_0[4748]); 
    assign out[1319] = layer_0[7998] & ~layer_0[2105]; 
    assign out[1320] = layer_0[2668] & ~layer_0[653]; 
    assign out[1321] = layer_0[2346] ^ layer_0[2362]; 
    assign out[1322] = ~(layer_0[6976] ^ layer_0[4455]); 
    assign out[1323] = ~(layer_0[5434] ^ layer_0[5924]); 
    assign out[1324] = ~layer_0[4409]; 
    assign out[1325] = ~(layer_0[1921] ^ layer_0[3482]); 
    assign out[1326] = layer_0[1220] ^ layer_0[462]; 
    assign out[1327] = layer_0[2228] ^ layer_0[367]; 
    assign out[1328] = ~(layer_0[2525] ^ layer_0[1675]); 
    assign out[1329] = layer_0[4323] ^ layer_0[6891]; 
    assign out[1330] = layer_0[6860] ^ layer_0[455]; 
    assign out[1331] = ~(layer_0[6132] ^ layer_0[4500]); 
    assign out[1332] = ~layer_0[4203] | (layer_0[1455] & layer_0[4203]); 
    assign out[1333] = layer_0[3069] & layer_0[382]; 
    assign out[1334] = layer_0[2525] & layer_0[6451]; 
    assign out[1335] = layer_0[3245] | layer_0[1390]; 
    assign out[1336] = ~layer_0[5094]; 
    assign out[1337] = layer_0[7894] ^ layer_0[6388]; 
    assign out[1338] = layer_0[4991] | layer_0[3594]; 
    assign out[1339] = ~(layer_0[5861] ^ layer_0[4702]); 
    assign out[1340] = layer_0[365]; 
    assign out[1341] = layer_0[6879] ^ layer_0[6936]; 
    assign out[1342] = ~(layer_0[2175] ^ layer_0[3635]); 
    assign out[1343] = layer_0[6441] ^ layer_0[2595]; 
    assign out[1344] = layer_0[5114] ^ layer_0[353]; 
    assign out[1345] = ~(layer_0[3297] | layer_0[2791]); 
    assign out[1346] = ~layer_0[2684]; 
    assign out[1347] = layer_0[3320] ^ layer_0[2358]; 
    assign out[1348] = layer_0[7312] ^ layer_0[7749]; 
    assign out[1349] = layer_0[2496] & ~layer_0[6696]; 
    assign out[1350] = ~(layer_0[1334] ^ layer_0[4316]); 
    assign out[1351] = ~layer_0[6774]; 
    assign out[1352] = ~layer_0[7962] | (layer_0[7962] & layer_0[925]); 
    assign out[1353] = layer_0[2503] ^ layer_0[4091]; 
    assign out[1354] = layer_0[345] ^ layer_0[3276]; 
    assign out[1355] = ~(layer_0[4216] ^ layer_0[2974]); 
    assign out[1356] = ~(layer_0[3193] ^ layer_0[4817]); 
    assign out[1357] = ~layer_0[1773]; 
    assign out[1358] = layer_0[3588] ^ layer_0[6669]; 
    assign out[1359] = layer_0[6288] ^ layer_0[7566]; 
    assign out[1360] = ~(layer_0[7001] ^ layer_0[6749]); 
    assign out[1361] = ~(layer_0[4888] ^ layer_0[4632]); 
    assign out[1362] = layer_0[4928]; 
    assign out[1363] = ~(layer_0[7329] | layer_0[4223]); 
    assign out[1364] = layer_0[1450]; 
    assign out[1365] = ~layer_0[7759] | (layer_0[5464] & layer_0[7759]); 
    assign out[1366] = layer_0[3579]; 
    assign out[1367] = ~(layer_0[6151] | layer_0[6815]); 
    assign out[1368] = ~layer_0[7010] | (layer_0[7010] & layer_0[3708]); 
    assign out[1369] = layer_0[2263] ^ layer_0[5845]; 
    assign out[1370] = ~layer_0[6536]; 
    assign out[1371] = ~(layer_0[2509] ^ layer_0[2099]); 
    assign out[1372] = layer_0[5173]; 
    assign out[1373] = layer_0[1837] | layer_0[5900]; 
    assign out[1374] = ~(layer_0[2551] ^ layer_0[6874]); 
    assign out[1375] = layer_0[5818] ^ layer_0[6328]; 
    assign out[1376] = layer_0[6179] & ~layer_0[4483]; 
    assign out[1377] = layer_0[4584] & layer_0[1223]; 
    assign out[1378] = layer_0[7442] ^ layer_0[5553]; 
    assign out[1379] = ~layer_0[2865]; 
    assign out[1380] = layer_0[2029] ^ layer_0[509]; 
    assign out[1381] = ~(layer_0[988] ^ layer_0[6087]); 
    assign out[1382] = layer_0[1054] & ~layer_0[530]; 
    assign out[1383] = ~layer_0[5996] | (layer_0[3971] & layer_0[5996]); 
    assign out[1384] = layer_0[3724] & ~layer_0[4596]; 
    assign out[1385] = layer_0[4179] ^ layer_0[4445]; 
    assign out[1386] = layer_0[6530]; 
    assign out[1387] = layer_0[6572] ^ layer_0[4684]; 
    assign out[1388] = layer_0[6300]; 
    assign out[1389] = layer_0[7984] & ~layer_0[852]; 
    assign out[1390] = ~layer_0[4833]; 
    assign out[1391] = layer_0[3840] ^ layer_0[5604]; 
    assign out[1392] = layer_0[1021] ^ layer_0[4102]; 
    assign out[1393] = ~layer_0[3415] | (layer_0[6179] & layer_0[3415]); 
    assign out[1394] = ~layer_0[4902]; 
    assign out[1395] = layer_0[920] & ~layer_0[5465]; 
    assign out[1396] = layer_0[5110] & ~layer_0[2949]; 
    assign out[1397] = ~layer_0[1507]; 
    assign out[1398] = ~(layer_0[1518] | layer_0[3531]); 
    assign out[1399] = ~(layer_0[5780] & layer_0[2726]); 
    assign out[1400] = ~layer_0[2671]; 
    assign out[1401] = ~layer_0[7703]; 
    assign out[1402] = layer_0[3477] & layer_0[5846]; 
    assign out[1403] = ~(layer_0[6214] ^ layer_0[7284]); 
    assign out[1404] = ~(layer_0[7297] ^ layer_0[7470]); 
    assign out[1405] = layer_0[6456] ^ layer_0[1805]; 
    assign out[1406] = layer_0[2006] ^ layer_0[6935]; 
    assign out[1407] = ~(layer_0[2366] | layer_0[1863]); 
    assign out[1408] = layer_0[6027] ^ layer_0[6589]; 
    assign out[1409] = ~(layer_0[2466] ^ layer_0[4243]); 
    assign out[1410] = layer_0[337] & ~layer_0[6268]; 
    assign out[1411] = layer_0[7408] ^ layer_0[6281]; 
    assign out[1412] = ~(layer_0[7101] ^ layer_0[4746]); 
    assign out[1413] = layer_0[531] ^ layer_0[5927]; 
    assign out[1414] = layer_0[4898] ^ layer_0[4680]; 
    assign out[1415] = layer_0[305] ^ layer_0[6069]; 
    assign out[1416] = layer_0[2999] & layer_0[6375]; 
    assign out[1417] = layer_0[6029] & layer_0[6933]; 
    assign out[1418] = layer_0[7450] ^ layer_0[1024]; 
    assign out[1419] = ~layer_0[4569] | (layer_0[1467] & layer_0[4569]); 
    assign out[1420] = ~(layer_0[7793] ^ layer_0[3895]); 
    assign out[1421] = layer_0[4118] & ~layer_0[7462]; 
    assign out[1422] = ~(layer_0[778] | layer_0[5428]); 
    assign out[1423] = ~(layer_0[7006] ^ layer_0[7537]); 
    assign out[1424] = layer_0[5585] | layer_0[4292]; 
    assign out[1425] = layer_0[2097]; 
    assign out[1426] = ~(layer_0[2189] ^ layer_0[3367]); 
    assign out[1427] = layer_0[529] & layer_0[71]; 
    assign out[1428] = ~(layer_0[182] | layer_0[5935]); 
    assign out[1429] = ~(layer_0[5683] ^ layer_0[977]); 
    assign out[1430] = ~layer_0[586] | (layer_0[586] & layer_0[2004]); 
    assign out[1431] = ~(layer_0[6950] ^ layer_0[4100]); 
    assign out[1432] = layer_0[7701]; 
    assign out[1433] = layer_0[7555] ^ layer_0[5988]; 
    assign out[1434] = ~layer_0[6606]; 
    assign out[1435] = ~(layer_0[6783] ^ layer_0[1670]); 
    assign out[1436] = layer_0[585] ^ layer_0[934]; 
    assign out[1437] = layer_0[5150] & layer_0[1855]; 
    assign out[1438] = layer_0[7923] ^ layer_0[974]; 
    assign out[1439] = ~layer_0[4004] | (layer_0[4004] & layer_0[4869]); 
    assign out[1440] = layer_0[162] ^ layer_0[3121]; 
    assign out[1441] = layer_0[3855] & ~layer_0[5012]; 
    assign out[1442] = layer_0[5825] ^ layer_0[158]; 
    assign out[1443] = ~layer_0[3959] | (layer_0[4104] & layer_0[3959]); 
    assign out[1444] = layer_0[7015] | layer_0[2618]; 
    assign out[1445] = ~(layer_0[1543] ^ layer_0[1333]); 
    assign out[1446] = ~(layer_0[2541] ^ layer_0[2691]); 
    assign out[1447] = layer_0[3209] & layer_0[2340]; 
    assign out[1448] = layer_0[3339] ^ layer_0[4728]; 
    assign out[1449] = layer_0[7402] ^ layer_0[2978]; 
    assign out[1450] = ~(layer_0[3135] ^ layer_0[880]); 
    assign out[1451] = ~(layer_0[1289] ^ layer_0[6797]); 
    assign out[1452] = ~layer_0[2886]; 
    assign out[1453] = ~(layer_0[1644] ^ layer_0[865]); 
    assign out[1454] = ~(layer_0[3182] & layer_0[458]); 
    assign out[1455] = layer_0[5692] ^ layer_0[2944]; 
    assign out[1456] = ~(layer_0[4439] & layer_0[5038]); 
    assign out[1457] = ~(layer_0[4241] ^ layer_0[7633]); 
    assign out[1458] = ~(layer_0[6349] | layer_0[4317]); 
    assign out[1459] = ~layer_0[2353] | (layer_0[2353] & layer_0[3788]); 
    assign out[1460] = layer_0[2542] ^ layer_0[2707]; 
    assign out[1461] = ~layer_0[4519]; 
    assign out[1462] = ~(layer_0[3442] ^ layer_0[7755]); 
    assign out[1463] = layer_0[6442] & layer_0[891]; 
    assign out[1464] = ~(layer_0[6912] ^ layer_0[3287]); 
    assign out[1465] = ~layer_0[1743] | (layer_0[4977] & layer_0[1743]); 
    assign out[1466] = layer_0[3919] ^ layer_0[6465]; 
    assign out[1467] = ~(layer_0[7049] ^ layer_0[5034]); 
    assign out[1468] = ~(layer_0[1547] ^ layer_0[7826]); 
    assign out[1469] = ~(layer_0[4670] & layer_0[5293]); 
    assign out[1470] = layer_0[290] & ~layer_0[1749]; 
    assign out[1471] = layer_0[5558] ^ layer_0[1920]; 
    assign out[1472] = ~layer_0[4711] | (layer_0[705] & layer_0[4711]); 
    assign out[1473] = ~(layer_0[3021] ^ layer_0[2165]); 
    assign out[1474] = ~(layer_0[4520] ^ layer_0[3372]); 
    assign out[1475] = layer_0[149]; 
    assign out[1476] = layer_0[3172] ^ layer_0[2380]; 
    assign out[1477] = layer_0[6750] ^ layer_0[961]; 
    assign out[1478] = layer_0[6360]; 
    assign out[1479] = ~(layer_0[2799] ^ layer_0[624]); 
    assign out[1480] = layer_0[6329]; 
    assign out[1481] = layer_0[591]; 
    assign out[1482] = layer_0[7873] ^ layer_0[2598]; 
    assign out[1483] = ~(layer_0[4757] ^ layer_0[2108]); 
    assign out[1484] = ~(layer_0[7746] | layer_0[7187]); 
    assign out[1485] = layer_0[7003] & ~layer_0[7456]; 
    assign out[1486] = ~(layer_0[273] ^ layer_0[7841]); 
    assign out[1487] = layer_0[2081] & layer_0[1054]; 
    assign out[1488] = layer_0[2430] ^ layer_0[2834]; 
    assign out[1489] = layer_0[4776] ^ layer_0[4302]; 
    assign out[1490] = ~(layer_0[2980] ^ layer_0[336]); 
    assign out[1491] = ~(layer_0[7126] ^ layer_0[2356]); 
    assign out[1492] = ~layer_0[3852]; 
    assign out[1493] = layer_0[751]; 
    assign out[1494] = ~(layer_0[5653] & layer_0[4899]); 
    assign out[1495] = layer_0[5137] ^ layer_0[6244]; 
    assign out[1496] = layer_0[6245] & ~layer_0[4533]; 
    assign out[1497] = ~layer_0[5493]; 
    assign out[1498] = ~layer_0[5562] | (layer_0[2946] & layer_0[5562]); 
    assign out[1499] = layer_0[7733] | layer_0[3618]; 
    assign out[1500] = layer_0[1272]; 
    assign out[1501] = layer_0[481]; 
    assign out[1502] = ~(layer_0[1483] | layer_0[4378]); 
    assign out[1503] = ~(layer_0[5383] & layer_0[5514]); 
    assign out[1504] = layer_0[4816] ^ layer_0[5714]; 
    assign out[1505] = layer_0[2027] ^ layer_0[4278]; 
    assign out[1506] = ~(layer_0[7202] ^ layer_0[4129]); 
    assign out[1507] = ~(layer_0[2532] & layer_0[2955]); 
    assign out[1508] = layer_0[7414] ^ layer_0[4877]; 
    assign out[1509] = ~(layer_0[2276] ^ layer_0[4726]); 
    assign out[1510] = layer_0[2627] | layer_0[4499]; 
    assign out[1511] = layer_0[817] & ~layer_0[7575]; 
    assign out[1512] = layer_0[3803] & layer_0[4956]; 
    assign out[1513] = layer_0[4254] | layer_0[5926]; 
    assign out[1514] = layer_0[3674] & layer_0[508]; 
    assign out[1515] = layer_0[7279] ^ layer_0[7549]; 
    assign out[1516] = layer_0[4086] ^ layer_0[5555]; 
    assign out[1517] = ~layer_0[4335]; 
    assign out[1518] = layer_0[1757]; 
    assign out[1519] = ~layer_0[6232]; 
    assign out[1520] = layer_0[6337] & ~layer_0[3029]; 
    assign out[1521] = layer_0[588] ^ layer_0[4148]; 
    assign out[1522] = ~layer_0[3344]; 
    assign out[1523] = ~layer_0[1597] | (layer_0[6147] & layer_0[1597]); 
    assign out[1524] = ~(layer_0[4795] | layer_0[5348]); 
    assign out[1525] = ~(layer_0[1318] | layer_0[3524]); 
    assign out[1526] = layer_0[7931] & ~layer_0[6926]; 
    assign out[1527] = ~(layer_0[7878] ^ layer_0[2586]); 
    assign out[1528] = layer_0[4261] & layer_0[6516]; 
    assign out[1529] = layer_0[631] & ~layer_0[6991]; 
    assign out[1530] = ~(layer_0[1899] ^ layer_0[4038]); 
    assign out[1531] = layer_0[2918]; 
    assign out[1532] = ~layer_0[6027]; 
    assign out[1533] = layer_0[3587]; 
    assign out[1534] = layer_0[2762] & ~layer_0[7274]; 
    assign out[1535] = ~layer_0[3159]; 
    assign out[1536] = layer_0[6450] & layer_0[3056]; 
    assign out[1537] = ~(layer_0[287] ^ layer_0[2313]); 
    assign out[1538] = ~(layer_0[747] ^ layer_0[2114]); 
    assign out[1539] = layer_0[3644] ^ layer_0[1248]; 
    assign out[1540] = layer_0[6056] & layer_0[4793]; 
    assign out[1541] = layer_0[7730] & ~layer_0[4810]; 
    assign out[1542] = layer_0[3888]; 
    assign out[1543] = layer_0[753]; 
    assign out[1544] = ~layer_0[874] | (layer_0[4261] & layer_0[874]); 
    assign out[1545] = layer_0[3570] ^ layer_0[2917]; 
    assign out[1546] = layer_0[5642]; 
    assign out[1547] = ~(layer_0[1697] & layer_0[6162]); 
    assign out[1548] = ~(layer_0[5949] ^ layer_0[2423]); 
    assign out[1549] = ~(layer_0[2975] | layer_0[1299]); 
    assign out[1550] = ~(layer_0[1865] ^ layer_0[359]); 
    assign out[1551] = layer_0[5997] ^ layer_0[6420]; 
    assign out[1552] = ~(layer_0[1348] ^ layer_0[5105]); 
    assign out[1553] = ~(layer_0[2237] ^ layer_0[1553]); 
    assign out[1554] = layer_0[7750] ^ layer_0[5177]; 
    assign out[1555] = ~(layer_0[6518] ^ layer_0[3691]); 
    assign out[1556] = layer_0[7040]; 
    assign out[1557] = ~(layer_0[5398] ^ layer_0[4022]); 
    assign out[1558] = layer_0[4205] ^ layer_0[3740]; 
    assign out[1559] = ~(layer_0[3939] ^ layer_0[6765]); 
    assign out[1560] = ~(layer_0[1022] & layer_0[390]); 
    assign out[1561] = layer_0[2538] ^ layer_0[7266]; 
    assign out[1562] = ~(layer_0[2741] ^ layer_0[2122]); 
    assign out[1563] = ~(layer_0[7359] ^ layer_0[1956]); 
    assign out[1564] = ~layer_0[7724]; 
    assign out[1565] = ~layer_0[7035]; 
    assign out[1566] = layer_0[6419] | layer_0[7962]; 
    assign out[1567] = layer_0[35] & ~layer_0[1178]; 
    assign out[1568] = layer_0[3019] ^ layer_0[3144]; 
    assign out[1569] = ~(layer_0[2631] & layer_0[1312]); 
    assign out[1570] = ~(layer_0[620] ^ layer_0[5443]); 
    assign out[1571] = ~(layer_0[4068] ^ layer_0[5656]); 
    assign out[1572] = layer_0[1924] ^ layer_0[332]; 
    assign out[1573] = layer_0[864]; 
    assign out[1574] = layer_0[6457] ^ layer_0[2388]; 
    assign out[1575] = layer_0[2814] & ~layer_0[6522]; 
    assign out[1576] = layer_0[1804] | layer_0[1120]; 
    assign out[1577] = ~(layer_0[5729] & layer_0[1218]); 
    assign out[1578] = layer_0[2197] ^ layer_0[933]; 
    assign out[1579] = ~(layer_0[5139] ^ layer_0[6105]); 
    assign out[1580] = ~(layer_0[672] | layer_0[2749]); 
    assign out[1581] = ~layer_0[5877] | (layer_0[5877] & layer_0[6845]); 
    assign out[1582] = layer_0[134]; 
    assign out[1583] = layer_0[54]; 
    assign out[1584] = ~layer_0[5228]; 
    assign out[1585] = ~(layer_0[7855] ^ layer_0[5166]); 
    assign out[1586] = layer_0[1409] ^ layer_0[6823]; 
    assign out[1587] = ~layer_0[473] | (layer_0[5089] & layer_0[473]); 
    assign out[1588] = ~(layer_0[1986] ^ layer_0[1187]); 
    assign out[1589] = layer_0[2261] ^ layer_0[3216]; 
    assign out[1590] = layer_0[5570] ^ layer_0[6969]; 
    assign out[1591] = layer_0[6325]; 
    assign out[1592] = layer_0[4067] ^ layer_0[519]; 
    assign out[1593] = layer_0[3173]; 
    assign out[1594] = layer_0[4371] ^ layer_0[3843]; 
    assign out[1595] = ~(layer_0[1815] | layer_0[3715]); 
    assign out[1596] = ~(layer_0[2734] ^ layer_0[4054]); 
    assign out[1597] = layer_0[3014] & layer_0[7615]; 
    assign out[1598] = layer_0[4627] ^ layer_0[4058]; 
    assign out[1599] = layer_0[3951] & ~layer_0[4782]; 
    assign out[1600] = layer_0[7486]; 
    assign out[1601] = layer_0[1843]; 
    assign out[1602] = layer_0[3883] & layer_0[2535]; 
    assign out[1603] = layer_0[1267]; 
    assign out[1604] = ~(layer_0[6965] | layer_0[3118]); 
    assign out[1605] = ~(layer_0[2317] ^ layer_0[2032]); 
    assign out[1606] = layer_0[5764]; 
    assign out[1607] = layer_0[5384] ^ layer_0[45]; 
    assign out[1608] = layer_0[3162] ^ layer_0[1188]; 
    assign out[1609] = layer_0[1050] & ~layer_0[3039]; 
    assign out[1610] = layer_0[6407]; 
    assign out[1611] = ~(layer_0[2853] ^ layer_0[2740]); 
    assign out[1612] = ~layer_0[2558]; 
    assign out[1613] = ~layer_0[3370]; 
    assign out[1614] = ~(layer_0[5160] & layer_0[4035]); 
    assign out[1615] = layer_0[5799]; 
    assign out[1616] = layer_0[921]; 
    assign out[1617] = layer_0[6924] & layer_0[5805]; 
    assign out[1618] = ~(layer_0[693] & layer_0[6295]); 
    assign out[1619] = layer_0[2005] & ~layer_0[1147]; 
    assign out[1620] = ~(layer_0[3185] & layer_0[2123]); 
    assign out[1621] = layer_0[7361] ^ layer_0[776]; 
    assign out[1622] = ~layer_0[4821] | (layer_0[4821] & layer_0[495]); 
    assign out[1623] = ~layer_0[843]; 
    assign out[1624] = layer_0[7679] & layer_0[7443]; 
    assign out[1625] = ~(layer_0[2588] & layer_0[5668]); 
    assign out[1626] = layer_0[6505] & ~layer_0[2816]; 
    assign out[1627] = ~layer_0[5280] | (layer_0[2873] & layer_0[5280]); 
    assign out[1628] = ~(layer_0[4603] ^ layer_0[5913]); 
    assign out[1629] = layer_0[6273]; 
    assign out[1630] = ~(layer_0[5132] ^ layer_0[4059]); 
    assign out[1631] = ~layer_0[566] | (layer_0[5503] & layer_0[566]); 
    assign out[1632] = ~(layer_0[6023] | layer_0[7769]); 
    assign out[1633] = ~layer_0[6046]; 
    assign out[1634] = layer_0[1438] & layer_0[5902]; 
    assign out[1635] = layer_0[4511]; 
    assign out[1636] = layer_0[3662] ^ layer_0[6234]; 
    assign out[1637] = layer_0[5751] & ~layer_0[3162]; 
    assign out[1638] = ~(layer_0[6066] | layer_0[5136]); 
    assign out[1639] = layer_0[4681] ^ layer_0[3934]; 
    assign out[1640] = ~layer_0[7356]; 
    assign out[1641] = layer_0[599]; 
    assign out[1642] = ~(layer_0[6393] ^ layer_0[6706]); 
    assign out[1643] = layer_0[3989] | layer_0[1871]; 
    assign out[1644] = layer_0[4605] ^ layer_0[1141]; 
    assign out[1645] = ~(layer_0[5356] ^ layer_0[3417]); 
    assign out[1646] = ~(layer_0[6893] ^ layer_0[4631]); 
    assign out[1647] = ~(layer_0[245] ^ layer_0[2989]); 
    assign out[1648] = ~layer_0[1113] | (layer_0[1113] & layer_0[6386]); 
    assign out[1649] = layer_0[5591] | layer_0[5579]; 
    assign out[1650] = layer_0[7905] & layer_0[1475]; 
    assign out[1651] = layer_0[1138] ^ layer_0[6384]; 
    assign out[1652] = ~layer_0[6635]; 
    assign out[1653] = layer_0[900] ^ layer_0[5126]; 
    assign out[1654] = layer_0[2753] ^ layer_0[1925]; 
    assign out[1655] = ~layer_0[1071] | (layer_0[6742] & layer_0[1071]); 
    assign out[1656] = ~(layer_0[4373] ^ layer_0[206]); 
    assign out[1657] = ~(layer_0[2534] & layer_0[3730]); 
    assign out[1658] = ~layer_0[7205]; 
    assign out[1659] = layer_0[802] ^ layer_0[7183]; 
    assign out[1660] = ~(layer_0[3772] ^ layer_0[914]); 
    assign out[1661] = ~(layer_0[3453] ^ layer_0[3249]); 
    assign out[1662] = ~layer_0[2907]; 
    assign out[1663] = layer_0[7277] & ~layer_0[4139]; 
    assign out[1664] = ~(layer_0[6977] ^ layer_0[2800]); 
    assign out[1665] = ~layer_0[4217]; 
    assign out[1666] = layer_0[2682] | layer_0[3036]; 
    assign out[1667] = ~layer_0[451]; 
    assign out[1668] = ~layer_0[2736] | (layer_0[2736] & layer_0[1765]); 
    assign out[1669] = layer_0[7525] ^ layer_0[1648]; 
    assign out[1670] = ~(layer_0[5068] ^ layer_0[3125]); 
    assign out[1671] = layer_0[2098] ^ layer_0[949]; 
    assign out[1672] = layer_0[6835]; 
    assign out[1673] = layer_0[4393] & ~layer_0[6971]; 
    assign out[1674] = ~(layer_0[3984] ^ layer_0[853]); 
    assign out[1675] = layer_0[5071]; 
    assign out[1676] = ~(layer_0[7867] | layer_0[2446]); 
    assign out[1677] = ~layer_0[4349]; 
    assign out[1678] = layer_0[2636]; 
    assign out[1679] = layer_0[1469] ^ layer_0[1061]; 
    assign out[1680] = ~(layer_0[4597] ^ layer_0[6452]); 
    assign out[1681] = ~(layer_0[3830] ^ layer_0[3983]); 
    assign out[1682] = ~(layer_0[207] ^ layer_0[4534]); 
    assign out[1683] = ~(layer_0[3593] ^ layer_0[6461]); 
    assign out[1684] = layer_0[2648]; 
    assign out[1685] = ~layer_0[3157]; 
    assign out[1686] = ~layer_0[2336]; 
    assign out[1687] = ~layer_0[7350] | (layer_0[1699] & layer_0[7350]); 
    assign out[1688] = ~(layer_0[4230] ^ layer_0[2985]); 
    assign out[1689] = layer_0[4743]; 
    assign out[1690] = ~(layer_0[7229] ^ layer_0[343]); 
    assign out[1691] = ~layer_0[3041]; 
    assign out[1692] = ~(layer_0[3122] ^ layer_0[2339]); 
    assign out[1693] = ~(layer_0[3236] ^ layer_0[6313]); 
    assign out[1694] = ~layer_0[1368] | (layer_0[7093] & layer_0[1368]); 
    assign out[1695] = ~(layer_0[7422] ^ layer_0[4604]); 
    assign out[1696] = layer_0[2311]; 
    assign out[1697] = ~(layer_0[1681] ^ layer_0[4109]); 
    assign out[1698] = layer_0[6590] ^ layer_0[2036]; 
    assign out[1699] = ~(layer_0[5987] | layer_0[6309]); 
    assign out[1700] = ~layer_0[6623] | (layer_0[5525] & layer_0[6623]); 
    assign out[1701] = layer_0[2935] & ~layer_0[5943]; 
    assign out[1702] = ~layer_0[854] | (layer_0[854] & layer_0[2370]); 
    assign out[1703] = ~(layer_0[2773] ^ layer_0[2795]); 
    assign out[1704] = layer_0[285]; 
    assign out[1705] = ~(layer_0[2925] ^ layer_0[967]); 
    assign out[1706] = ~(layer_0[5119] ^ layer_0[6396]); 
    assign out[1707] = ~layer_0[3062] | (layer_0[3521] & layer_0[3062]); 
    assign out[1708] = layer_0[2823] ^ layer_0[4187]; 
    assign out[1709] = ~layer_0[2050] | (layer_0[4930] & layer_0[2050]); 
    assign out[1710] = ~(layer_0[138] ^ layer_0[5932]); 
    assign out[1711] = ~layer_0[6509] | (layer_0[361] & layer_0[6509]); 
    assign out[1712] = layer_0[4015] ^ layer_0[6987]; 
    assign out[1713] = layer_0[2286] & ~layer_0[4011]; 
    assign out[1714] = ~layer_0[3516] | (layer_0[3516] & layer_0[6277]); 
    assign out[1715] = layer_0[4130]; 
    assign out[1716] = layer_0[2890] ^ layer_0[2955]; 
    assign out[1717] = layer_0[4224] ^ layer_0[5240]; 
    assign out[1718] = layer_0[1769] ^ layer_0[642]; 
    assign out[1719] = layer_0[7669] ^ layer_0[5668]; 
    assign out[1720] = layer_0[7547] ^ layer_0[7657]; 
    assign out[1721] = ~(layer_0[3528] ^ layer_0[7772]); 
    assign out[1722] = layer_0[7933] | layer_0[3342]; 
    assign out[1723] = ~layer_0[5622]; 
    assign out[1724] = ~(layer_0[5135] ^ layer_0[4353]); 
    assign out[1725] = ~(layer_0[4221] ^ layer_0[5772]); 
    assign out[1726] = layer_0[1840] ^ layer_0[7940]; 
    assign out[1727] = ~layer_0[2939] | (layer_0[6671] & layer_0[2939]); 
    assign out[1728] = layer_0[3101] ^ layer_0[7481]; 
    assign out[1729] = layer_0[1969] | layer_0[2757]; 
    assign out[1730] = layer_0[4886] & ~layer_0[7140]; 
    assign out[1731] = layer_0[3884]; 
    assign out[1732] = layer_0[1950] & layer_0[72]; 
    assign out[1733] = ~layer_0[3568] | (layer_0[4334] & layer_0[3568]); 
    assign out[1734] = ~(layer_0[7254] ^ layer_0[772]); 
    assign out[1735] = ~(layer_0[7804] ^ layer_0[1152]); 
    assign out[1736] = layer_0[234]; 
    assign out[1737] = layer_0[923] ^ layer_0[4906]; 
    assign out[1738] = layer_0[1616] ^ layer_0[5096]; 
    assign out[1739] = ~(layer_0[1937] ^ layer_0[7839]); 
    assign out[1740] = layer_0[4551]; 
    assign out[1741] = ~layer_0[5874] | (layer_0[5955] & layer_0[5874]); 
    assign out[1742] = ~(layer_0[7215] & layer_0[5046]); 
    assign out[1743] = ~(layer_0[4151] ^ layer_0[71]); 
    assign out[1744] = layer_0[3404] & layer_0[896]; 
    assign out[1745] = ~(layer_0[6169] ^ layer_0[7549]); 
    assign out[1746] = layer_0[1149] | layer_0[3680]; 
    assign out[1747] = ~(layer_0[6339] ^ layer_0[7454]); 
    assign out[1748] = ~(layer_0[7458] | layer_0[4653]); 
    assign out[1749] = layer_0[4938]; 
    assign out[1750] = layer_0[1706] ^ layer_0[2304]; 
    assign out[1751] = layer_0[2283]; 
    assign out[1752] = layer_0[3124]; 
    assign out[1753] = layer_0[3200] ^ layer_0[6901]; 
    assign out[1754] = ~(layer_0[1223] ^ layer_0[1309]); 
    assign out[1755] = layer_0[3777] ^ layer_0[3096]; 
    assign out[1756] = ~(layer_0[3597] ^ layer_0[7323]); 
    assign out[1757] = ~layer_0[5021]; 
    assign out[1758] = layer_0[2518] ^ layer_0[5770]; 
    assign out[1759] = layer_0[2244] & layer_0[1981]; 
    assign out[1760] = ~(layer_0[5964] ^ layer_0[5485]); 
    assign out[1761] = layer_0[7531]; 
    assign out[1762] = layer_0[2244]; 
    assign out[1763] = ~(layer_0[666] | layer_0[3086]); 
    assign out[1764] = layer_0[5317] & ~layer_0[2998]; 
    assign out[1765] = ~(layer_0[139] ^ layer_0[2976]); 
    assign out[1766] = ~(layer_0[1901] ^ layer_0[7489]); 
    assign out[1767] = layer_0[1803] ^ layer_0[1949]; 
    assign out[1768] = layer_0[3749]; 
    assign out[1769] = ~layer_0[2950] | (layer_0[2950] & layer_0[121]); 
    assign out[1770] = ~(layer_0[5269] ^ layer_0[4623]); 
    assign out[1771] = ~(layer_0[1852] & layer_0[2802]); 
    assign out[1772] = ~layer_0[2343]; 
    assign out[1773] = ~(layer_0[6743] ^ layer_0[4233]); 
    assign out[1774] = layer_0[3310] & ~layer_0[6592]; 
    assign out[1775] = ~layer_0[2809]; 
    assign out[1776] = ~(layer_0[5801] ^ layer_0[4483]); 
    assign out[1777] = ~(layer_0[4546] ^ layer_0[5021]); 
    assign out[1778] = ~(layer_0[5895] ^ layer_0[438]); 
    assign out[1779] = ~layer_0[420]; 
    assign out[1780] = layer_0[5679]; 
    assign out[1781] = layer_0[6588]; 
    assign out[1782] = ~layer_0[4238]; 
    assign out[1783] = ~(layer_0[2157] ^ layer_0[4571]); 
    assign out[1784] = layer_0[3352] ^ layer_0[1996]; 
    assign out[1785] = ~(layer_0[6044] ^ layer_0[5557]); 
    assign out[1786] = layer_0[3914] & ~layer_0[666]; 
    assign out[1787] = ~(layer_0[1521] ^ layer_0[535]); 
    assign out[1788] = ~layer_0[7145] | (layer_0[7145] & layer_0[4481]); 
    assign out[1789] = ~layer_0[5381] | (layer_0[7740] & layer_0[5381]); 
    assign out[1790] = ~(layer_0[7097] ^ layer_0[1774]); 
    assign out[1791] = ~(layer_0[6683] ^ layer_0[6641]); 
    assign out[1792] = ~(layer_0[7967] ^ layer_0[1062]); 
    assign out[1793] = layer_0[7716] & ~layer_0[4365]; 
    assign out[1794] = ~layer_0[6954] | (layer_0[6954] & layer_0[7561]); 
    assign out[1795] = layer_0[2416] ^ layer_0[7135]; 
    assign out[1796] = layer_0[3957]; 
    assign out[1797] = layer_0[2564] | layer_0[7983]; 
    assign out[1798] = ~(layer_0[5797] ^ layer_0[2187]); 
    assign out[1799] = layer_0[6979] & ~layer_0[3379]; 
    assign out[1800] = layer_0[6195]; 
    assign out[1801] = layer_0[1034] ^ layer_0[7301]; 
    assign out[1802] = ~layer_0[5610] | (layer_0[5610] & layer_0[3924]); 
    assign out[1803] = layer_0[3591] & layer_0[6977]; 
    assign out[1804] = ~(layer_0[304] ^ layer_0[5331]); 
    assign out[1805] = ~(layer_0[5044] ^ layer_0[7416]); 
    assign out[1806] = layer_0[4874] ^ layer_0[2199]; 
    assign out[1807] = ~layer_0[4843] | (layer_0[4843] & layer_0[5073]); 
    assign out[1808] = ~(layer_0[5186] ^ layer_0[7853]); 
    assign out[1809] = ~(layer_0[7971] ^ layer_0[2232]); 
    assign out[1810] = layer_0[5257]; 
    assign out[1811] = layer_0[3419] & layer_0[4280]; 
    assign out[1812] = ~layer_0[23] | (layer_0[23] & layer_0[5644]); 
    assign out[1813] = ~(layer_0[5174] ^ layer_0[2878]); 
    assign out[1814] = layer_0[4014] & ~layer_0[6096]; 
    assign out[1815] = layer_0[151] & layer_0[6745]; 
    assign out[1816] = layer_0[554] ^ layer_0[7114]; 
    assign out[1817] = layer_0[4176]; 
    assign out[1818] = layer_0[1479] ^ layer_0[2365]; 
    assign out[1819] = layer_0[4701]; 
    assign out[1820] = layer_0[7216] ^ layer_0[1282]; 
    assign out[1821] = layer_0[4031]; 
    assign out[1822] = layer_0[5092] ^ layer_0[2500]; 
    assign out[1823] = layer_0[7178] ^ layer_0[924]; 
    assign out[1824] = layer_0[5598]; 
    assign out[1825] = layer_0[737] ^ layer_0[4929]; 
    assign out[1826] = ~layer_0[6646]; 
    assign out[1827] = layer_0[7095] ^ layer_0[4469]; 
    assign out[1828] = ~(layer_0[5651] ^ layer_0[5446]); 
    assign out[1829] = ~layer_0[5115] | (layer_0[4907] & layer_0[5115]); 
    assign out[1830] = layer_0[324]; 
    assign out[1831] = layer_0[4988] ^ layer_0[2888]; 
    assign out[1832] = ~layer_0[3350] | (layer_0[3350] & layer_0[6779]); 
    assign out[1833] = ~layer_0[5014] | (layer_0[5271] & layer_0[5014]); 
    assign out[1834] = ~layer_0[2375]; 
    assign out[1835] = ~(layer_0[5791] | layer_0[5276]); 
    assign out[1836] = ~layer_0[2692] | (layer_0[2692] & layer_0[3657]); 
    assign out[1837] = layer_0[6065]; 
    assign out[1838] = layer_0[4411] & ~layer_0[4139]; 
    assign out[1839] = layer_0[4548] ^ layer_0[3008]; 
    assign out[1840] = layer_0[756] ^ layer_0[4984]; 
    assign out[1841] = ~(layer_0[395] ^ layer_0[6975]); 
    assign out[1842] = ~(layer_0[2973] & layer_0[5388]); 
    assign out[1843] = ~(layer_0[949] ^ layer_0[2956]); 
    assign out[1844] = ~layer_0[2856] | (layer_0[5587] & layer_0[2856]); 
    assign out[1845] = layer_0[7786] & ~layer_0[4440]; 
    assign out[1846] = layer_0[3530] ^ layer_0[4084]; 
    assign out[1847] = ~(layer_0[1057] ^ layer_0[4040]); 
    assign out[1848] = ~layer_0[7532]; 
    assign out[1849] = ~(layer_0[5203] & layer_0[775]); 
    assign out[1850] = ~(layer_0[5182] & layer_0[1903]); 
    assign out[1851] = ~layer_0[3355]; 
    assign out[1852] = layer_0[5248]; 
    assign out[1853] = layer_0[4882] & layer_0[7768]; 
    assign out[1854] = layer_0[2352] & ~layer_0[907]; 
    assign out[1855] = ~(layer_0[6032] ^ layer_0[6409]); 
    assign out[1856] = layer_0[4725] ^ layer_0[6180]; 
    assign out[1857] = layer_0[1668]; 
    assign out[1858] = layer_0[4404]; 
    assign out[1859] = layer_0[5113] & ~layer_0[5080]; 
    assign out[1860] = ~(layer_0[7117] | layer_0[7169]); 
    assign out[1861] = layer_0[3987] ^ layer_0[6793]; 
    assign out[1862] = layer_0[1417] & ~layer_0[6916]; 
    assign out[1863] = layer_0[6031] & layer_0[7357]; 
    assign out[1864] = ~(layer_0[1174] ^ layer_0[232]); 
    assign out[1865] = layer_0[4802] ^ layer_0[6447]; 
    assign out[1866] = layer_0[2125]; 
    assign out[1867] = layer_0[3147] & layer_0[5917]; 
    assign out[1868] = ~(layer_0[978] ^ layer_0[4521]); 
    assign out[1869] = ~layer_0[157]; 
    assign out[1870] = layer_0[4004] ^ layer_0[3892]; 
    assign out[1871] = ~(layer_0[6492] ^ layer_0[1165]); 
    assign out[1872] = layer_0[4535] ^ layer_0[4143]; 
    assign out[1873] = layer_0[2064] ^ layer_0[642]; 
    assign out[1874] = ~(layer_0[3188] ^ layer_0[2789]); 
    assign out[1875] = layer_0[5631]; 
    assign out[1876] = ~(layer_0[3997] ^ layer_0[4252]); 
    assign out[1877] = layer_0[4573] & ~layer_0[7263]; 
    assign out[1878] = layer_0[1185] ^ layer_0[7758]; 
    assign out[1879] = layer_0[2487] & ~layer_0[4574]; 
    assign out[1880] = ~(layer_0[1000] ^ layer_0[3301]); 
    assign out[1881] = ~layer_0[6587] | (layer_0[4978] & layer_0[6587]); 
    assign out[1882] = ~layer_0[4279] | (layer_0[2803] & layer_0[4279]); 
    assign out[1883] = layer_0[7397] ^ layer_0[756]; 
    assign out[1884] = layer_0[4295] ^ layer_0[7428]; 
    assign out[1885] = ~(layer_0[4457] & layer_0[315]); 
    assign out[1886] = layer_0[7988] & ~layer_0[81]; 
    assign out[1887] = layer_0[1148] & ~layer_0[1661]; 
    assign out[1888] = layer_0[4996] ^ layer_0[1674]; 
    assign out[1889] = ~(layer_0[7431] ^ layer_0[5775]); 
    assign out[1890] = ~(layer_0[4942] ^ layer_0[6447]); 
    assign out[1891] = ~layer_0[1105]; 
    assign out[1892] = ~layer_0[4430]; 
    assign out[1893] = ~(layer_0[5255] ^ layer_0[7773]); 
    assign out[1894] = layer_0[3483] | layer_0[1842]; 
    assign out[1895] = layer_0[7581] ^ layer_0[6547]; 
    assign out[1896] = ~(layer_0[1979] | layer_0[3865]); 
    assign out[1897] = layer_0[3374]; 
    assign out[1898] = ~(layer_0[6135] ^ layer_0[4363]); 
    assign out[1899] = ~layer_0[4310]; 
    assign out[1900] = layer_0[7112] & layer_0[7778]; 
    assign out[1901] = layer_0[4405] ^ layer_0[3384]; 
    assign out[1902] = ~layer_0[7150]; 
    assign out[1903] = ~(layer_0[2896] ^ layer_0[1628]); 
    assign out[1904] = layer_0[2041] ^ layer_0[2086]; 
    assign out[1905] = layer_0[4985]; 
    assign out[1906] = ~layer_0[441]; 
    assign out[1907] = layer_0[2170] ^ layer_0[6512]; 
    assign out[1908] = ~(layer_0[1715] ^ layer_0[5457]); 
    assign out[1909] = layer_0[1661]; 
    assign out[1910] = ~(layer_0[1376] ^ layer_0[2512]); 
    assign out[1911] = layer_0[4621] | layer_0[32]; 
    assign out[1912] = layer_0[5490]; 
    assign out[1913] = layer_0[4944]; 
    assign out[1914] = ~layer_0[3052] | (layer_0[3052] & layer_0[5870]); 
    assign out[1915] = ~(layer_0[6653] | layer_0[4801]); 
    assign out[1916] = layer_0[1995]; 
    assign out[1917] = layer_0[2961] ^ layer_0[1519]; 
    assign out[1918] = layer_0[4134] ^ layer_0[3165]; 
    assign out[1919] = ~(layer_0[5757] ^ layer_0[1183]); 
    assign out[1920] = layer_0[935] ^ layer_0[590]; 
    assign out[1921] = ~layer_0[1735] | (layer_0[3752] & layer_0[1735]); 
    assign out[1922] = ~(layer_0[1443] ^ layer_0[2402]); 
    assign out[1923] = layer_0[5284] ^ layer_0[6590]; 
    assign out[1924] = layer_0[2324] | layer_0[6679]; 
    assign out[1925] = ~layer_0[1041]; 
    assign out[1926] = layer_0[1926]; 
    assign out[1927] = ~layer_0[5011]; 
    assign out[1928] = layer_0[735] ^ layer_0[1572]; 
    assign out[1929] = layer_0[6812] ^ layer_0[568]; 
    assign out[1930] = layer_0[393] ^ layer_0[1831]; 
    assign out[1931] = ~(layer_0[7811] | layer_0[3683]); 
    assign out[1932] = ~(layer_0[719] ^ layer_0[5936]); 
    assign out[1933] = ~(layer_0[7579] | layer_0[6271]); 
    assign out[1934] = ~layer_0[5814]; 
    assign out[1935] = layer_0[7937] | layer_0[5886]; 
    assign out[1936] = layer_0[6085] & ~layer_0[5430]; 
    assign out[1937] = layer_0[3560] | layer_0[5457]; 
    assign out[1938] = ~(layer_0[208] ^ layer_0[4366]); 
    assign out[1939] = ~(layer_0[7909] & layer_0[5651]); 
    assign out[1940] = ~(layer_0[137] ^ layer_0[6225]); 
    assign out[1941] = layer_0[1420] | layer_0[4021]; 
    assign out[1942] = layer_0[5610] ^ layer_0[5573]; 
    assign out[1943] = ~(layer_0[1202] & layer_0[3693]); 
    assign out[1944] = ~(layer_0[3831] | layer_0[3758]); 
    assign out[1945] = ~layer_0[46] | (layer_0[46] & layer_0[6806]); 
    assign out[1946] = ~(layer_0[92] ^ layer_0[2143]); 
    assign out[1947] = layer_0[675]; 
    assign out[1948] = ~(layer_0[3108] ^ layer_0[3185]); 
    assign out[1949] = layer_0[1516] ^ layer_0[7948]; 
    assign out[1950] = layer_0[214] ^ layer_0[598]; 
    assign out[1951] = ~layer_0[2342]; 
    assign out[1952] = ~layer_0[6008]; 
    assign out[1953] = layer_0[5586] & ~layer_0[5471]; 
    assign out[1954] = layer_0[790] & layer_0[4289]; 
    assign out[1955] = layer_0[5447] & layer_0[6700]; 
    assign out[1956] = layer_0[6290] ^ layer_0[912]; 
    assign out[1957] = ~(layer_0[4155] ^ layer_0[5635]); 
    assign out[1958] = layer_0[4663] & ~layer_0[6665]; 
    assign out[1959] = layer_0[3266] ^ layer_0[6276]; 
    assign out[1960] = ~(layer_0[764] ^ layer_0[7117]); 
    assign out[1961] = ~layer_0[394] | (layer_0[2037] & layer_0[394]); 
    assign out[1962] = layer_0[5962]; 
    assign out[1963] = layer_0[6249] & ~layer_0[1111]; 
    assign out[1964] = layer_0[6507]; 
    assign out[1965] = ~layer_0[4250]; 
    assign out[1966] = ~layer_0[3999] | (layer_0[7478] & layer_0[3999]); 
    assign out[1967] = ~(layer_0[755] | layer_0[2909]); 
    assign out[1968] = ~(layer_0[1565] & layer_0[7781]); 
    assign out[1969] = layer_0[2847] & layer_0[3440]; 
    assign out[1970] = ~(layer_0[4606] ^ layer_0[6175]); 
    assign out[1971] = ~layer_0[1167] | (layer_0[1167] & layer_0[757]); 
    assign out[1972] = ~layer_0[5401] | (layer_0[5401] & layer_0[6934]); 
    assign out[1973] = layer_0[1784] ^ layer_0[2453]; 
    assign out[1974] = ~layer_0[4912] | (layer_0[154] & layer_0[4912]); 
    assign out[1975] = layer_0[1817] & layer_0[5290]; 
    assign out[1976] = layer_0[4852] ^ layer_0[4703]; 
    assign out[1977] = ~(layer_0[6607] & layer_0[4331]); 
    assign out[1978] = ~(layer_0[3853] ^ layer_0[827]); 
    assign out[1979] = ~layer_0[6882] | (layer_0[6882] & layer_0[2628]); 
    assign out[1980] = layer_0[3183] ^ layer_0[66]; 
    assign out[1981] = layer_0[6964] & ~layer_0[7827]; 
    assign out[1982] = layer_0[3226] ^ layer_0[1357]; 
    assign out[1983] = layer_0[3763] ^ layer_0[662]; 
    assign out[1984] = layer_0[6150] & layer_0[5040]; 
    assign out[1985] = ~(layer_0[1136] ^ layer_0[6012]); 
    assign out[1986] = layer_0[4489] ^ layer_0[5852]; 
    assign out[1987] = ~(layer_0[4128] ^ layer_0[3198]); 
    assign out[1988] = layer_0[4956] ^ layer_0[7750]; 
    assign out[1989] = layer_0[5312] & ~layer_0[647]; 
    assign out[1990] = ~(layer_0[2456] ^ layer_0[3905]); 
    assign out[1991] = ~layer_0[6854] | (layer_0[6854] & layer_0[1475]); 
    assign out[1992] = ~(layer_0[5620] ^ layer_0[1642]); 
    assign out[1993] = layer_0[6028] ^ layer_0[2894]; 
    assign out[1994] = layer_0[2158] ^ layer_0[2977]; 
    assign out[1995] = ~(layer_0[3928] ^ layer_0[467]); 
    assign out[1996] = layer_0[2321] & layer_0[1005]; 
    assign out[1997] = ~(layer_0[3314] ^ layer_0[5973]); 
    assign out[1998] = ~layer_0[4773] | (layer_0[4773] & layer_0[7175]); 
    assign out[1999] = layer_0[3553] ^ layer_0[1152]; 
    assign out[2000] = ~layer_0[10] | (layer_0[10] & layer_0[3443]); 
    assign out[2001] = layer_0[1109]; 
    assign out[2002] = ~(layer_0[4980] ^ layer_0[152]); 
    assign out[2003] = ~(layer_0[6142] ^ layer_0[667]); 
    assign out[2004] = layer_0[6617] ^ layer_0[837]; 
    assign out[2005] = ~(layer_0[1478] | layer_0[7276]); 
    assign out[2006] = layer_0[3402] ^ layer_0[5049]; 
    assign out[2007] = ~(layer_0[5595] ^ layer_0[3262]); 
    assign out[2008] = ~(layer_0[4502] ^ layer_0[4518]); 
    assign out[2009] = layer_0[364] ^ layer_0[6458]; 
    assign out[2010] = ~(layer_0[2412] ^ layer_0[7649]); 
    assign out[2011] = layer_0[699]; 
    assign out[2012] = layer_0[4187] ^ layer_0[3629]; 
    assign out[2013] = ~(layer_0[7702] ^ layer_0[4857]); 
    assign out[2014] = ~(layer_0[62] ^ layer_0[1915]); 
    assign out[2015] = ~(layer_0[7853] & layer_0[1351]); 
    assign out[2016] = ~layer_0[5349] | (layer_0[5349] & layer_0[3352]); 
    assign out[2017] = ~layer_0[805]; 
    assign out[2018] = layer_0[7753] ^ layer_0[1695]; 
    assign out[2019] = ~(layer_0[3369] ^ layer_0[810]); 
    assign out[2020] = ~(layer_0[2259] & layer_0[3455]); 
    assign out[2021] = layer_0[1073] | layer_0[1671]; 
    assign out[2022] = layer_0[4174] | layer_0[6482]; 
    assign out[2023] = ~layer_0[2719]; 
    assign out[2024] = layer_0[2704] | layer_0[543]; 
    assign out[2025] = layer_0[2174] ^ layer_0[1429]; 
    assign out[2026] = ~(layer_0[5057] ^ layer_0[379]); 
    assign out[2027] = layer_0[6462]; 
    assign out[2028] = ~(layer_0[6460] ^ layer_0[5342]); 
    assign out[2029] = ~(layer_0[4157] | layer_0[3090]); 
    assign out[2030] = layer_0[4403]; 
    assign out[2031] = layer_0[5551] ^ layer_0[3240]; 
    assign out[2032] = ~(layer_0[6776] | layer_0[6601]); 
    assign out[2033] = ~layer_0[2681] | (layer_0[4338] & layer_0[2681]); 
    assign out[2034] = layer_0[875]; 
    assign out[2035] = ~(layer_0[1994] & layer_0[2660]); 
    assign out[2036] = 1'b1; 
    assign out[2037] = layer_0[6909]; 
    assign out[2038] = layer_0[674] ^ layer_0[1633]; 
    assign out[2039] = layer_0[237] | layer_0[1750]; 
    assign out[2040] = ~layer_0[4273] | (layer_0[4273] & layer_0[6174]); 
    assign out[2041] = ~(layer_0[4402] & layer_0[1182]); 
    assign out[2042] = ~(layer_0[443] ^ layer_0[2335]); 
    assign out[2043] = layer_0[5536] & ~layer_0[742]; 
    assign out[2044] = layer_0[7147] ^ layer_0[3615]; 
    assign out[2045] = ~(layer_0[943] ^ layer_0[664]); 
    assign out[2046] = ~(layer_0[6114] ^ layer_0[1930]); 
    assign out[2047] = layer_0[5896] & ~layer_0[7982]; 
    assign out[2048] = layer_0[5346] ^ layer_0[3032]; 
    assign out[2049] = ~(layer_0[27] | layer_0[6294]); 
    assign out[2050] = layer_0[3564] ^ layer_0[3726]; 
    assign out[2051] = ~(layer_0[3787] ^ layer_0[1582]); 
    assign out[2052] = ~(layer_0[3672] | layer_0[6785]); 
    assign out[2053] = layer_0[1180] ^ layer_0[6167]; 
    assign out[2054] = layer_0[7786] ^ layer_0[1946]; 
    assign out[2055] = layer_0[3329]; 
    assign out[2056] = layer_0[521]; 
    assign out[2057] = 1'b0; 
    assign out[2058] = ~layer_0[5792]; 
    assign out[2059] = layer_0[6449] & layer_0[6152]; 
    assign out[2060] = layer_0[1788] & ~layer_0[6928]; 
    assign out[2061] = layer_0[7515] & ~layer_0[6492]; 
    assign out[2062] = layer_0[4736] ^ layer_0[6259]; 
    assign out[2063] = layer_0[3722] | layer_0[1252]; 
    assign out[2064] = layer_0[6881] | layer_0[5193]; 
    assign out[2065] = ~layer_0[7829]; 
    assign out[2066] = layer_0[18] ^ layer_0[4712]; 
    assign out[2067] = layer_0[987] & ~layer_0[1815]; 
    assign out[2068] = ~(layer_0[1444] ^ layer_0[426]); 
    assign out[2069] = layer_0[1982] ^ layer_0[509]; 
    assign out[2070] = ~(layer_0[1696] ^ layer_0[723]); 
    assign out[2071] = layer_0[926] ^ layer_0[7967]; 
    assign out[2072] = ~(layer_0[5170] ^ layer_0[4910]); 
    assign out[2073] = layer_0[1825] ^ layer_0[1756]; 
    assign out[2074] = ~(layer_0[501] ^ layer_0[5267]); 
    assign out[2075] = ~(layer_0[6754] | layer_0[3407]); 
    assign out[2076] = layer_0[1171] & layer_0[4042]; 
    assign out[2077] = ~(layer_0[5803] | layer_0[4622]); 
    assign out[2078] = ~(layer_0[6956] ^ layer_0[1608]); 
    assign out[2079] = ~(layer_0[2954] ^ layer_0[6681]); 
    assign out[2080] = layer_0[7847] ^ layer_0[2226]; 
    assign out[2081] = layer_0[7433] & ~layer_0[3239]; 
    assign out[2082] = ~layer_0[3815]; 
    assign out[2083] = ~(layer_0[1857] ^ layer_0[5728]); 
    assign out[2084] = layer_0[4198]; 
    assign out[2085] = layer_0[3291] & ~layer_0[7595]; 
    assign out[2086] = 1'b0; 
    assign out[2087] = ~(layer_0[4876] ^ layer_0[391]); 
    assign out[2088] = ~(layer_0[2281] ^ layer_0[7735]); 
    assign out[2089] = layer_0[2505] & ~layer_0[2264]; 
    assign out[2090] = ~(layer_0[3060] ^ layer_0[1408]); 
    assign out[2091] = layer_0[4608] ^ layer_0[5199]; 
    assign out[2092] = ~layer_0[378]; 
    assign out[2093] = layer_0[6241] ^ layer_0[4895]; 
    assign out[2094] = layer_0[6168] & ~layer_0[1888]; 
    assign out[2095] = ~(layer_0[1973] ^ layer_0[5978]); 
    assign out[2096] = ~layer_0[2031]; 
    assign out[2097] = ~(layer_0[6377] | layer_0[3214]); 
    assign out[2098] = layer_0[4431] ^ layer_0[2806]; 
    assign out[2099] = layer_0[979]; 
    assign out[2100] = layer_0[5602] & layer_0[7590]; 
    assign out[2101] = layer_0[6762] ^ layer_0[7360]; 
    assign out[2102] = ~layer_0[3935] | (layer_0[3935] & layer_0[3356]); 
    assign out[2103] = layer_0[2750] ^ layer_0[1255]; 
    assign out[2104] = layer_0[747] ^ layer_0[1238]; 
    assign out[2105] = layer_0[663] & ~layer_0[5299]; 
    assign out[2106] = layer_0[6809] & ~layer_0[2610]; 
    assign out[2107] = layer_0[6138] ^ layer_0[5067]; 
    assign out[2108] = layer_0[2779] & ~layer_0[5619]; 
    assign out[2109] = layer_0[5866] & ~layer_0[4456]; 
    assign out[2110] = ~layer_0[4436]; 
    assign out[2111] = layer_0[6123] ^ layer_0[3122]; 
    assign out[2112] = ~(layer_0[7717] ^ layer_0[7522]); 
    assign out[2113] = ~(layer_0[2347] | layer_0[1153]); 
    assign out[2114] = layer_0[3046] ^ layer_0[2821]; 
    assign out[2115] = layer_0[1453] & layer_0[4962]; 
    assign out[2116] = ~layer_0[148]; 
    assign out[2117] = ~(layer_0[6048] | layer_0[6308]); 
    assign out[2118] = layer_0[911] & ~layer_0[6915]; 
    assign out[2119] = layer_0[6960] ^ layer_0[7827]; 
    assign out[2120] = layer_0[6812] | layer_0[4704]; 
    assign out[2121] = ~(layer_0[1923] ^ layer_0[968]); 
    assign out[2122] = layer_0[1976] | layer_0[1907]; 
    assign out[2123] = layer_0[5687] ^ layer_0[3388]; 
    assign out[2124] = ~(layer_0[6407] ^ layer_0[4017]); 
    assign out[2125] = ~(layer_0[4760] ^ layer_0[1999]); 
    assign out[2126] = layer_0[2701] & ~layer_0[6081]; 
    assign out[2127] = layer_0[3143] ^ layer_0[6380]; 
    assign out[2128] = layer_0[7015]; 
    assign out[2129] = layer_0[3216] ^ layer_0[1945]; 
    assign out[2130] = ~layer_0[1567]; 
    assign out[2131] = ~(layer_0[2497] ^ layer_0[3510]); 
    assign out[2132] = layer_0[2267] ^ layer_0[1256]; 
    assign out[2133] = layer_0[6353] ^ layer_0[7380]; 
    assign out[2134] = ~layer_0[5822]; 
    assign out[2135] = ~(layer_0[7146] ^ layer_0[704]); 
    assign out[2136] = layer_0[3773] ^ layer_0[6929]; 
    assign out[2137] = ~layer_0[4565]; 
    assign out[2138] = layer_0[6698] | layer_0[3945]; 
    assign out[2139] = layer_0[2109] | layer_0[5977]; 
    assign out[2140] = ~layer_0[3716] | (layer_0[3716] & layer_0[4675]); 
    assign out[2141] = ~(layer_0[1238] ^ layer_0[6636]); 
    assign out[2142] = ~layer_0[5975]; 
    assign out[2143] = ~layer_0[1827]; 
    assign out[2144] = ~(layer_0[2259] & layer_0[2907]); 
    assign out[2145] = layer_0[2895] ^ layer_0[6553]; 
    assign out[2146] = layer_0[3257] & layer_0[3327]; 
    assign out[2147] = ~(layer_0[3962] | layer_0[702]); 
    assign out[2148] = layer_0[5167] ^ layer_0[6770]; 
    assign out[2149] = layer_0[5649]; 
    assign out[2150] = layer_0[1602] ^ layer_0[5013]; 
    assign out[2151] = ~layer_0[7904] | (layer_0[5158] & layer_0[7904]); 
    assign out[2152] = ~(layer_0[6158] | layer_0[6838]); 
    assign out[2153] = layer_0[3175]; 
    assign out[2154] = layer_0[2822] & ~layer_0[4169]; 
    assign out[2155] = layer_0[3582] & ~layer_0[497]; 
    assign out[2156] = ~(layer_0[1410] ^ layer_0[5624]); 
    assign out[2157] = ~layer_0[6331]; 
    assign out[2158] = layer_0[2020]; 
    assign out[2159] = layer_0[1150] ^ layer_0[75]; 
    assign out[2160] = layer_0[6322] & ~layer_0[700]; 
    assign out[2161] = layer_0[5221] & layer_0[7972]; 
    assign out[2162] = layer_0[1792] & ~layer_0[5010]; 
    assign out[2163] = ~(layer_0[7401] ^ layer_0[5390]); 
    assign out[2164] = layer_0[6299] & ~layer_0[5056]; 
    assign out[2165] = layer_0[2060] ^ layer_0[6491]; 
    assign out[2166] = layer_0[673] & ~layer_0[3793]; 
    assign out[2167] = ~(layer_0[6171] ^ layer_0[498]); 
    assign out[2168] = layer_0[3900] & ~layer_0[2869]; 
    assign out[2169] = layer_0[6648] ^ layer_0[1]; 
    assign out[2170] = layer_0[5029] ^ layer_0[5801]; 
    assign out[2171] = layer_0[5058] ^ layer_0[4797]; 
    assign out[2172] = layer_0[3849]; 
    assign out[2173] = layer_0[5242] ^ layer_0[5350]; 
    assign out[2174] = layer_0[2151] ^ layer_0[7761]; 
    assign out[2175] = ~(layer_0[1400] | layer_0[2476]); 
    assign out[2176] = layer_0[2536]; 
    assign out[2177] = ~(layer_0[4196] ^ layer_0[1155]); 
    assign out[2178] = layer_0[4023] & layer_0[5810]; 
    assign out[2179] = ~(layer_0[27] ^ layer_0[2969]); 
    assign out[2180] = ~(layer_0[3982] ^ layer_0[1573]); 
    assign out[2181] = ~(layer_0[228] ^ layer_0[2417]); 
    assign out[2182] = ~(layer_0[1195] ^ layer_0[3105]); 
    assign out[2183] = layer_0[3269] ^ layer_0[5202]; 
    assign out[2184] = ~(layer_0[6643] & layer_0[3712]); 
    assign out[2185] = layer_0[4172] ^ layer_0[2811]; 
    assign out[2186] = layer_0[288] & ~layer_0[5046]; 
    assign out[2187] = layer_0[215] & ~layer_0[5081]; 
    assign out[2188] = ~layer_0[7118] | (layer_0[7118] & layer_0[4445]); 
    assign out[2189] = 1'b1; 
    assign out[2190] = layer_0[5443] ^ layer_0[302]; 
    assign out[2191] = layer_0[2536] ^ layer_0[1226]; 
    assign out[2192] = ~(layer_0[4027] ^ layer_0[796]); 
    assign out[2193] = ~layer_0[2807]; 
    assign out[2194] = layer_0[6066] & ~layer_0[5495]; 
    assign out[2195] = layer_0[1848] & ~layer_0[3345]; 
    assign out[2196] = layer_0[6178] & ~layer_0[4123]; 
    assign out[2197] = ~(layer_0[197] ^ layer_0[2158]); 
    assign out[2198] = layer_0[7704] & ~layer_0[3611]; 
    assign out[2199] = ~(layer_0[1659] ^ layer_0[490]); 
    assign out[2200] = ~(layer_0[4066] & layer_0[7460]); 
    assign out[2201] = layer_0[6850]; 
    assign out[2202] = layer_0[119] ^ layer_0[4572]; 
    assign out[2203] = layer_0[4853]; 
    assign out[2204] = ~(layer_0[3634] ^ layer_0[4528]); 
    assign out[2205] = ~(layer_0[5728] ^ layer_0[6469]); 
    assign out[2206] = ~(layer_0[3048] | layer_0[6836]); 
    assign out[2207] = layer_0[7048]; 
    assign out[2208] = layer_0[6568] | layer_0[4764]; 
    assign out[2209] = ~(layer_0[842] ^ layer_0[1927]); 
    assign out[2210] = layer_0[7783] ^ layer_0[4140]; 
    assign out[2211] = layer_0[1070] | layer_0[352]; 
    assign out[2212] = ~(layer_0[7123] ^ layer_0[1729]); 
    assign out[2213] = layer_0[3291] & ~layer_0[6122]; 
    assign out[2214] = layer_0[2771] & layer_0[3484]; 
    assign out[2215] = layer_0[6310] & layer_0[4003]; 
    assign out[2216] = ~(layer_0[1812] ^ layer_0[4189]); 
    assign out[2217] = layer_0[6230] ^ layer_0[1554]; 
    assign out[2218] = ~(layer_0[3195] | layer_0[1896]); 
    assign out[2219] = layer_0[264]; 
    assign out[2220] = ~layer_0[3707] | (layer_0[703] & layer_0[3707]); 
    assign out[2221] = layer_0[6921] ^ layer_0[3078]; 
    assign out[2222] = ~(layer_0[4880] ^ layer_0[6633]); 
    assign out[2223] = layer_0[7094] ^ layer_0[3656]; 
    assign out[2224] = layer_0[7138] ^ layer_0[1682]; 
    assign out[2225] = layer_0[1778] ^ layer_0[4870]; 
    assign out[2226] = ~(layer_0[4449] | layer_0[5008]); 
    assign out[2227] = layer_0[1799] ^ layer_0[5477]; 
    assign out[2228] = layer_0[3826] & layer_0[1687]; 
    assign out[2229] = ~layer_0[1440]; 
    assign out[2230] = ~layer_0[1491] | (layer_0[5655] & layer_0[1491]); 
    assign out[2231] = ~(layer_0[7390] ^ layer_0[4742]); 
    assign out[2232] = layer_0[698] ^ layer_0[6916]; 
    assign out[2233] = layer_0[3357] ^ layer_0[2902]; 
    assign out[2234] = layer_0[3972] ^ layer_0[3181]; 
    assign out[2235] = ~(layer_0[6670] ^ layer_0[4536]); 
    assign out[2236] = layer_0[7799] & ~layer_0[3094]; 
    assign out[2237] = ~layer_0[7250]; 
    assign out[2238] = layer_0[6269] & ~layer_0[2499]; 
    assign out[2239] = ~(layer_0[478] ^ layer_0[318]); 
    assign out[2240] = layer_0[316] & ~layer_0[6667]; 
    assign out[2241] = ~(layer_0[2133] ^ layer_0[5943]); 
    assign out[2242] = ~layer_0[1050] | (layer_0[5394] & layer_0[1050]); 
    assign out[2243] = layer_0[1213] ^ layer_0[4515]; 
    assign out[2244] = ~(layer_0[2530] ^ layer_0[372]); 
    assign out[2245] = ~(layer_0[7385] ^ layer_0[3083]); 
    assign out[2246] = ~layer_0[6829]; 
    assign out[2247] = layer_0[1609]; 
    assign out[2248] = ~layer_0[3689] | (layer_0[3689] & layer_0[7836]); 
    assign out[2249] = ~layer_0[4813]; 
    assign out[2250] = ~(layer_0[1944] ^ layer_0[1430]); 
    assign out[2251] = ~(layer_0[7090] ^ layer_0[4552]); 
    assign out[2252] = ~(layer_0[1121] ^ layer_0[2382]); 
    assign out[2253] = layer_0[5073] ^ layer_0[6112]; 
    assign out[2254] = layer_0[7156] ^ layer_0[3219]; 
    assign out[2255] = layer_0[6376] ^ layer_0[2562]; 
    assign out[2256] = ~layer_0[7303]; 
    assign out[2257] = layer_0[5067]; 
    assign out[2258] = layer_0[283]; 
    assign out[2259] = layer_0[2063]; 
    assign out[2260] = layer_0[2938] & ~layer_0[3462]; 
    assign out[2261] = layer_0[2072] & ~layer_0[386]; 
    assign out[2262] = ~layer_0[732] | (layer_0[406] & layer_0[732]); 
    assign out[2263] = ~layer_0[2840]; 
    assign out[2264] = ~(layer_0[1200] ^ layer_0[6137]); 
    assign out[2265] = layer_0[2597] ^ layer_0[5783]; 
    assign out[2266] = ~(layer_0[6370] ^ layer_0[7419]); 
    assign out[2267] = layer_0[6130]; 
    assign out[2268] = layer_0[5738] ^ layer_0[6084]; 
    assign out[2269] = ~layer_0[1093]; 
    assign out[2270] = ~(layer_0[2074] ^ layer_0[4584]); 
    assign out[2271] = layer_0[6183] ^ layer_0[937]; 
    assign out[2272] = ~(layer_0[6852] & layer_0[6788]); 
    assign out[2273] = ~(layer_0[7859] & layer_0[3158]); 
    assign out[2274] = layer_0[265] ^ layer_0[272]; 
    assign out[2275] = ~layer_0[7455] | (layer_0[7455] & layer_0[2584]); 
    assign out[2276] = ~layer_0[5487] | (layer_0[5487] & layer_0[2406]); 
    assign out[2277] = ~(layer_0[4778] ^ layer_0[4713]); 
    assign out[2278] = ~(layer_0[3192] ^ layer_0[3917]); 
    assign out[2279] = layer_0[4225] ^ layer_0[3052]; 
    assign out[2280] = ~layer_0[971]; 
    assign out[2281] = layer_0[2225] ^ layer_0[25]; 
    assign out[2282] = layer_0[4646] & layer_0[3231]; 
    assign out[2283] = layer_0[2870] ^ layer_0[6900]; 
    assign out[2284] = layer_0[7672] ^ layer_0[492]; 
    assign out[2285] = ~layer_0[1098]; 
    assign out[2286] = layer_0[6518] | layer_0[6724]; 
    assign out[2287] = layer_0[1910] ^ layer_0[4294]; 
    assign out[2288] = ~(layer_0[6701] ^ layer_0[3491]); 
    assign out[2289] = layer_0[7538] ^ layer_0[7236]; 
    assign out[2290] = ~(layer_0[4127] ^ layer_0[4741]); 
    assign out[2291] = ~(layer_0[4247] & layer_0[1746]); 
    assign out[2292] = layer_0[3366] ^ layer_0[2360]; 
    assign out[2293] = ~(layer_0[946] ^ layer_0[3496]); 
    assign out[2294] = layer_0[1556] & ~layer_0[2484]; 
    assign out[2295] = 1'b0; 
    assign out[2296] = ~(layer_0[1521] ^ layer_0[3546]); 
    assign out[2297] = ~(layer_0[4178] | layer_0[5759]); 
    assign out[2298] = layer_0[7584]; 
    assign out[2299] = ~(layer_0[354] ^ layer_0[2951]); 
    assign out[2300] = ~(layer_0[5521] ^ layer_0[258]); 
    assign out[2301] = ~layer_0[5184] | (layer_0[4963] & layer_0[5184]); 
    assign out[2302] = layer_0[1393]; 
    assign out[2303] = layer_0[3869] ^ layer_0[5441]; 
    assign out[2304] = ~(layer_0[5588] ^ layer_0[7288]); 
    assign out[2305] = ~(layer_0[1005] ^ layer_0[6666]); 
    assign out[2306] = layer_0[7951] ^ layer_0[276]; 
    assign out[2307] = ~(layer_0[2104] ^ layer_0[362]); 
    assign out[2308] = layer_0[6527] ^ layer_0[6133]; 
    assign out[2309] = ~(layer_0[4099] ^ layer_0[2367]); 
    assign out[2310] = layer_0[2619]; 
    assign out[2311] = ~(layer_0[5458] ^ layer_0[896]); 
    assign out[2312] = ~(layer_0[1834] ^ layer_0[6582]); 
    assign out[2313] = ~layer_0[5210]; 
    assign out[2314] = layer_0[4419] & ~layer_0[5899]; 
    assign out[2315] = layer_0[4274] & ~layer_0[363]; 
    assign out[2316] = ~(layer_0[3923] ^ layer_0[6768]); 
    assign out[2317] = ~layer_0[6306]; 
    assign out[2318] = layer_0[7545] & layer_0[789]; 
    assign out[2319] = layer_0[7812] & ~layer_0[4379]; 
    assign out[2320] = ~layer_0[2835]; 
    assign out[2321] = layer_0[3497] & ~layer_0[1456]; 
    assign out[2322] = layer_0[7333] & layer_0[3572]; 
    assign out[2323] = layer_0[1144] ^ layer_0[610]; 
    assign out[2324] = ~layer_0[752]; 
    assign out[2325] = ~(layer_0[1868] ^ layer_0[2964]); 
    assign out[2326] = layer_0[7663] ^ layer_0[2343]; 
    assign out[2327] = ~(layer_0[6802] ^ layer_0[6610]); 
    assign out[2328] = layer_0[2208] ^ layer_0[3618]; 
    assign out[2329] = ~(layer_0[5238] | layer_0[6064]); 
    assign out[2330] = ~layer_0[2065] | (layer_0[2065] & layer_0[1224]); 
    assign out[2331] = ~layer_0[3503] | (layer_0[7897] & layer_0[3503]); 
    assign out[2332] = layer_0[557]; 
    assign out[2333] = layer_0[4501] ^ layer_0[1623]; 
    assign out[2334] = layer_0[4268] & ~layer_0[61]; 
    assign out[2335] = ~layer_0[3405] | (layer_0[2045] & layer_0[3405]); 
    assign out[2336] = layer_0[7391] ^ layer_0[1754]; 
    assign out[2337] = 1'b1; 
    assign out[2338] = ~(layer_0[4530] & layer_0[4204]); 
    assign out[2339] = ~(layer_0[4701] ^ layer_0[4064]); 
    assign out[2340] = layer_0[2769] ^ layer_0[3513]; 
    assign out[2341] = layer_0[1311] ^ layer_0[5523]; 
    assign out[2342] = ~(layer_0[7665] | layer_0[194]); 
    assign out[2343] = layer_0[7993] ^ layer_0[6208]; 
    assign out[2344] = layer_0[965] & layer_0[4642]; 
    assign out[2345] = ~(layer_0[7204] ^ layer_0[696]); 
    assign out[2346] = layer_0[2459] ^ layer_0[2137]; 
    assign out[2347] = ~layer_0[795] | (layer_0[3227] & layer_0[795]); 
    assign out[2348] = ~(layer_0[3651] ^ layer_0[3387]); 
    assign out[2349] = ~layer_0[2922] | (layer_0[2922] & layer_0[5222]); 
    assign out[2350] = ~(layer_0[6955] & layer_0[1544]); 
    assign out[2351] = ~(layer_0[4762] ^ layer_0[2206]); 
    assign out[2352] = layer_0[3809] ^ layer_0[569]; 
    assign out[2353] = ~(layer_0[5104] ^ layer_0[7727]); 
    assign out[2354] = ~layer_0[5344]; 
    assign out[2355] = ~layer_0[5637]; 
    assign out[2356] = layer_0[5211] & layer_0[7530]; 
    assign out[2357] = layer_0[5734] & ~layer_0[4856]; 
    assign out[2358] = layer_0[6278] ^ layer_0[7369]; 
    assign out[2359] = layer_0[431] ^ layer_0[160]; 
    assign out[2360] = layer_0[7139] ^ layer_0[3397]; 
    assign out[2361] = ~(layer_0[2666] ^ layer_0[4214]); 
    assign out[2362] = ~layer_0[6332]; 
    assign out[2363] = layer_0[2864] & layer_0[3492]; 
    assign out[2364] = layer_0[633] | layer_0[2523]; 
    assign out[2365] = ~(layer_0[7311] ^ layer_0[5226]); 
    assign out[2366] = layer_0[547] ^ layer_0[1636]; 
    assign out[2367] = layer_0[6549] ^ layer_0[5872]; 
    assign out[2368] = layer_0[4664] & ~layer_0[4348]; 
    assign out[2369] = ~(layer_0[3343] ^ layer_0[1841]); 
    assign out[2370] = ~layer_0[4791] | (layer_0[7660] & layer_0[4791]); 
    assign out[2371] = layer_0[4346] & ~layer_0[6141]; 
    assign out[2372] = layer_0[731] | layer_0[3725]; 
    assign out[2373] = layer_0[7251] | layer_0[3138]; 
    assign out[2374] = layer_0[271] ^ layer_0[1529]; 
    assign out[2375] = layer_0[432] ^ layer_0[634]; 
    assign out[2376] = layer_0[4616] & layer_0[1605]; 
    assign out[2377] = layer_0[6103] & ~layer_0[4276]; 
    assign out[2378] = layer_0[4470] ^ layer_0[7079]; 
    assign out[2379] = layer_0[3265]; 
    assign out[2380] = ~layer_0[1362]; 
    assign out[2381] = layer_0[4024] & layer_0[3112]; 
    assign out[2382] = layer_0[7991] & layer_0[3894]; 
    assign out[2383] = ~layer_0[5524]; 
    assign out[2384] = layer_0[3823] ^ layer_0[3135]; 
    assign out[2385] = ~(layer_0[4472] ^ layer_0[6771]); 
    assign out[2386] = ~layer_0[2565] | (layer_0[835] & layer_0[2565]); 
    assign out[2387] = ~(layer_0[5403] ^ layer_0[4446]); 
    assign out[2388] = layer_0[4113]; 
    assign out[2389] = layer_0[4901] ^ layer_0[4339]; 
    assign out[2390] = layer_0[2404] ^ layer_0[3847]; 
    assign out[2391] = ~(layer_0[3903] | layer_0[2071]); 
    assign out[2392] = layer_0[4753]; 
    assign out[2393] = layer_0[6803] ^ layer_0[5432]; 
    assign out[2394] = layer_0[2567] ^ layer_0[6785]; 
    assign out[2395] = layer_0[7325] ^ layer_0[335]; 
    assign out[2396] = layer_0[7315] & ~layer_0[1643]; 
    assign out[2397] = layer_0[6586] & ~layer_0[7464]; 
    assign out[2398] = layer_0[2794] ^ layer_0[4505]; 
    assign out[2399] = layer_0[7300] ^ layer_0[285]; 
    assign out[2400] = layer_0[398] & layer_0[3064]; 
    assign out[2401] = ~(layer_0[3946] ^ layer_0[2144]); 
    assign out[2402] = layer_0[1386] & layer_0[303]; 
    assign out[2403] = ~(layer_0[3085] | layer_0[1592]); 
    assign out[2404] = layer_0[428] ^ layer_0[7176]; 
    assign out[2405] = layer_0[7020] ^ layer_0[7259]; 
    assign out[2406] = layer_0[69] & layer_0[4277]; 
    assign out[2407] = ~layer_0[1577]; 
    assign out[2408] = layer_0[3655] & ~layer_0[816]; 
    assign out[2409] = layer_0[4780]; 
    assign out[2410] = ~(layer_0[1414] | layer_0[7915]); 
    assign out[2411] = layer_0[6856] ^ layer_0[1775]; 
    assign out[2412] = layer_0[5106] ^ layer_0[5473]; 
    assign out[2413] = layer_0[7987] & ~layer_0[2290]; 
    assign out[2414] = layer_0[7526] ^ layer_0[1686]; 
    assign out[2415] = ~(layer_0[4210] & layer_0[6186]); 
    assign out[2416] = layer_0[4862] ^ layer_0[5613]; 
    assign out[2417] = layer_0[6559]; 
    assign out[2418] = ~layer_0[6369]; 
    assign out[2419] = layer_0[7774] ^ layer_0[3463]; 
    assign out[2420] = layer_0[6932] & layer_0[5582]; 
    assign out[2421] = layer_0[2216] & ~layer_0[652]; 
    assign out[2422] = ~(layer_0[7736] ^ layer_0[7033]); 
    assign out[2423] = ~(layer_0[4140] ^ layer_0[2010]); 
    assign out[2424] = layer_0[4453] ^ layer_0[1648]; 
    assign out[2425] = layer_0[4890] ^ layer_0[2612]; 
    assign out[2426] = ~(layer_0[7317] ^ layer_0[4184]); 
    assign out[2427] = ~(layer_0[2589] | layer_0[3391]); 
    assign out[2428] = layer_0[2566] & ~layer_0[4496]; 
    assign out[2429] = ~(layer_0[3156] | layer_0[3906]); 
    assign out[2430] = layer_0[2059]; 
    assign out[2431] = layer_0[3184] & layer_0[3836]; 
    assign out[2432] = layer_0[2480] ^ layer_0[208]; 
    assign out[2433] = layer_0[1613] ^ layer_0[6002]; 
    assign out[2434] = ~(layer_0[3452] ^ layer_0[3289]); 
    assign out[2435] = ~(layer_0[7133] ^ layer_0[7685]); 
    assign out[2436] = ~layer_0[6672]; 
    assign out[2437] = ~(layer_0[928] ^ layer_0[5367]); 
    assign out[2438] = ~layer_0[720] | (layer_0[720] & layer_0[7188]); 
    assign out[2439] = ~(layer_0[184] ^ layer_0[3602]); 
    assign out[2440] = layer_0[2540] & layer_0[5355]; 
    assign out[2441] = ~(layer_0[6846] ^ layer_0[4589]); 
    assign out[2442] = layer_0[546]; 
    assign out[2443] = ~layer_0[4761]; 
    assign out[2444] = ~(layer_0[2080] ^ layer_0[7491]); 
    assign out[2445] = ~(layer_0[1242] ^ layer_0[2805]); 
    assign out[2446] = layer_0[2555] ^ layer_0[5876]; 
    assign out[2447] = layer_0[1305] & layer_0[973]; 
    assign out[2448] = layer_0[7393] ^ layer_0[7200]; 
    assign out[2449] = layer_0[210] ^ layer_0[5377]; 
    assign out[2450] = layer_0[6257] ^ layer_0[7624]; 
    assign out[2451] = layer_0[578] & ~layer_0[4433]; 
    assign out[2452] = ~(layer_0[5100] ^ layer_0[3321]); 
    assign out[2453] = layer_0[3599] & layer_0[5724]; 
    assign out[2454] = layer_0[3457] ^ layer_0[1244]; 
    assign out[2455] = ~(layer_0[2227] ^ layer_0[6550]); 
    assign out[2456] = layer_0[2676] & ~layer_0[3292]; 
    assign out[2457] = layer_0[6842] ^ layer_0[5268]; 
    assign out[2458] = ~(layer_0[935] ^ layer_0[796]); 
    assign out[2459] = layer_0[3068] ^ layer_0[7077]; 
    assign out[2460] = layer_0[6514] & ~layer_0[4992]; 
    assign out[2461] = layer_0[5577] ^ layer_0[1304]; 
    assign out[2462] = layer_0[2424] & ~layer_0[606]; 
    assign out[2463] = layer_0[3766] ^ layer_0[4215]; 
    assign out[2464] = layer_0[6389] & layer_0[172]; 
    assign out[2465] = layer_0[7527] ^ layer_0[5320]; 
    assign out[2466] = layer_0[6165] ^ layer_0[7568]; 
    assign out[2467] = ~(layer_0[3664] & layer_0[1717]); 
    assign out[2468] = ~(layer_0[5762] & layer_0[6314]); 
    assign out[2469] = layer_0[4087] & ~layer_0[1669]; 
    assign out[2470] = ~layer_0[1708]; 
    assign out[2471] = layer_0[6775] ^ layer_0[5302]; 
    assign out[2472] = ~layer_0[7282]; 
    assign out[2473] = ~layer_0[1277] | (layer_0[1819] & layer_0[1277]); 
    assign out[2474] = ~(layer_0[5636] ^ layer_0[2873]); 
    assign out[2475] = layer_0[4671] ^ layer_0[1406]; 
    assign out[2476] = ~(layer_0[1125] ^ layer_0[4386]); 
    assign out[2477] = layer_0[4264] & ~layer_0[6875]; 
    assign out[2478] = ~(layer_0[291] ^ layer_0[5413]); 
    assign out[2479] = ~(layer_0[1097] ^ layer_0[6357]); 
    assign out[2480] = ~(layer_0[2728] ^ layer_0[1091]); 
    assign out[2481] = ~layer_0[3702]; 
    assign out[2482] = layer_0[6395] ^ layer_0[1207]; 
    assign out[2483] = ~(layer_0[5181] ^ layer_0[7852]); 
    assign out[2484] = ~(layer_0[7376] ^ layer_0[4396]); 
    assign out[2485] = layer_0[1531] & ~layer_0[6211]; 
    assign out[2486] = ~layer_0[7702]; 
    assign out[2487] = ~(layer_0[812] ^ layer_0[7264]); 
    assign out[2488] = layer_0[5520]; 
    assign out[2489] = layer_0[5632] ^ layer_0[4098]; 
    assign out[2490] = ~layer_0[6428] | (layer_0[6428] & layer_0[7447]); 
    assign out[2491] = ~(layer_0[798] ^ layer_0[4950]); 
    assign out[2492] = ~(layer_0[6343] ^ layer_0[1147]); 
    assign out[2493] = layer_0[7445]; 
    assign out[2494] = layer_0[2213] ^ layer_0[6970]; 
    assign out[2495] = ~(layer_0[3245] ^ layer_0[4056]); 
    assign out[2496] = ~layer_0[5440] | (layer_0[5512] & layer_0[5440]); 
    assign out[2497] = ~(layer_0[1874] ^ layer_0[5681]); 
    assign out[2498] = layer_0[6237] ^ layer_0[4916]; 
    assign out[2499] = ~layer_0[5534] | (layer_0[5534] & layer_0[7945]); 
    assign out[2500] = layer_0[1955] ^ layer_0[3263]; 
    assign out[2501] = layer_0[649] ^ layer_0[5499]; 
    assign out[2502] = layer_0[2718] ^ layer_0[4595]; 
    assign out[2503] = ~(layer_0[1796] ^ layer_0[499]); 
    assign out[2504] = layer_0[1359] | layer_0[356]; 
    assign out[2505] = ~(layer_0[417] ^ layer_0[2245]); 
    assign out[2506] = ~(layer_0[5047] ^ layer_0[5773]); 
    assign out[2507] = layer_0[7570] & ~layer_0[676]; 
    assign out[2508] = layer_0[645] | layer_0[5970]; 
    assign out[2509] = ~(layer_0[1425] & layer_0[1476]); 
    assign out[2510] = ~layer_0[3331] | (layer_0[7020] & layer_0[3331]); 
    assign out[2511] = layer_0[7187] ^ layer_0[3764]; 
    assign out[2512] = ~(layer_0[3805] ^ layer_0[3098]); 
    assign out[2513] = layer_0[6622] ^ layer_0[6573]; 
    assign out[2514] = layer_0[4918] ^ layer_0[5185]; 
    assign out[2515] = ~layer_0[4421] | (layer_0[4421] & layer_0[2547]); 
    assign out[2516] = layer_0[1677] ^ layer_0[6118]; 
    assign out[2517] = layer_0[7316] ^ layer_0[2514]; 
    assign out[2518] = ~(layer_0[6333] ^ layer_0[4447]); 
    assign out[2519] = ~(layer_0[4149] ^ layer_0[6695]); 
    assign out[2520] = layer_0[252] & layer_0[3779]; 
    assign out[2521] = layer_0[6481] & ~layer_0[5594]; 
    assign out[2522] = layer_0[1785] ^ layer_0[1542]; 
    assign out[2523] = ~layer_0[6684]; 
    assign out[2524] = layer_0[4036] ^ layer_0[3640]; 
    assign out[2525] = layer_0[3861] ^ layer_0[1413]; 
    assign out[2526] = ~layer_0[4390]; 
    assign out[2527] = layer_0[3983] ^ layer_0[4015]; 
    assign out[2528] = layer_0[4346] & layer_0[181]; 
    assign out[2529] = ~(layer_0[277] ^ layer_0[4153]); 
    assign out[2530] = ~layer_0[5322] | (layer_0[594] & layer_0[5322]); 
    assign out[2531] = ~(layer_0[1378] ^ layer_0[2456]); 
    assign out[2532] = layer_0[5059] ^ layer_0[1972]; 
    assign out[2533] = layer_0[2699] & ~layer_0[5286]; 
    assign out[2534] = layer_0[6093] ^ layer_0[6266]; 
    assign out[2535] = layer_0[7957]; 
    assign out[2536] = ~(layer_0[348] ^ layer_0[6070]); 
    assign out[2537] = layer_0[3991] ^ layer_0[4130]; 
    assign out[2538] = layer_0[5000]; 
    assign out[2539] = layer_0[4837] & ~layer_0[6647]; 
    assign out[2540] = ~(layer_0[5130] ^ layer_0[3869]); 
    assign out[2541] = layer_0[2185] ^ layer_0[5862]; 
    assign out[2542] = ~(layer_0[4572] | layer_0[7339]); 
    assign out[2543] = layer_0[2996] | layer_0[4559]; 
    assign out[2544] = layer_0[7344] & layer_0[239]; 
    assign out[2545] = layer_0[6582] ^ layer_0[3470]; 
    assign out[2546] = layer_0[7286] & ~layer_0[1489]; 
    assign out[2547] = ~layer_0[1702]; 
    assign out[2548] = layer_0[6034]; 
    assign out[2549] = layer_0[224] ^ layer_0[6942]; 
    assign out[2550] = layer_0[683] ^ layer_0[1711]; 
    assign out[2551] = ~(layer_0[1897] ^ layer_0[6145]); 
    assign out[2552] = layer_0[3306]; 
    assign out[2553] = ~layer_0[1968] | (layer_0[5516] & layer_0[1968]); 
    assign out[2554] = layer_0[1829] & layer_0[4488]; 
    assign out[2555] = ~(layer_0[1496] & layer_0[7025]); 
    assign out[2556] = layer_0[7406]; 
    assign out[2557] = ~layer_0[7821]; 
    assign out[2558] = ~layer_0[7050] | (layer_0[3890] & layer_0[7050]); 
    assign out[2559] = ~layer_0[2237] | (layer_0[7306] & layer_0[2237]); 
    assign out[2560] = layer_0[2546] & ~layer_0[7498]; 
    assign out[2561] = layer_0[541] ^ layer_0[4808]; 
    assign out[2562] = layer_0[745]; 
    assign out[2563] = ~layer_0[3099]; 
    assign out[2564] = layer_0[7238] ^ layer_0[5349]; 
    assign out[2565] = layer_0[6164]; 
    assign out[2566] = layer_0[6236] ^ layer_0[5370]; 
    assign out[2567] = layer_0[3066] | layer_0[1422]; 
    assign out[2568] = ~layer_0[2760]; 
    assign out[2569] = ~(layer_0[3323] ^ layer_0[6264]); 
    assign out[2570] = ~layer_0[6766] | (layer_0[6766] & layer_0[6242]); 
    assign out[2571] = layer_0[6862] ^ layer_0[641]; 
    assign out[2572] = ~(layer_0[6224] ^ layer_0[4047]); 
    assign out[2573] = ~layer_0[3170]; 
    assign out[2574] = layer_0[4162]; 
    assign out[2575] = layer_0[2217]; 
    assign out[2576] = ~layer_0[5375]; 
    assign out[2577] = layer_0[6082] & ~layer_0[2501]; 
    assign out[2578] = layer_0[6054] & layer_0[3992]; 
    assign out[2579] = ~layer_0[4] | (layer_0[3371] & layer_0[4]); 
    assign out[2580] = layer_0[1680] ^ layer_0[7116]; 
    assign out[2581] = layer_0[2209] & layer_0[4209]; 
    assign out[2582] = ~(layer_0[5356] & layer_0[2987]); 
    assign out[2583] = layer_0[2755] | layer_0[4838]; 
    assign out[2584] = ~layer_0[6159] | (layer_0[4006] & layer_0[6159]); 
    assign out[2585] = layer_0[3292]; 
    assign out[2586] = ~layer_0[670] | (layer_0[670] & layer_0[2602]); 
    assign out[2587] = layer_0[3807] | layer_0[5601]; 
    assign out[2588] = layer_0[2296] ^ layer_0[7543]; 
    assign out[2589] = layer_0[6194]; 
    assign out[2590] = layer_0[6118] & ~layer_0[5024]; 
    assign out[2591] = layer_0[3045] ^ layer_0[3822]; 
    assign out[2592] = layer_0[4479] ^ layer_0[6318]; 
    assign out[2593] = layer_0[1332] & layer_0[2225]; 
    assign out[2594] = layer_0[1689] ^ layer_0[5581]; 
    assign out[2595] = layer_0[1985] & ~layer_0[5289]; 
    assign out[2596] = ~(layer_0[536] ^ layer_0[4484]); 
    assign out[2597] = ~layer_0[439] | (layer_0[439] & layer_0[2011]); 
    assign out[2598] = layer_0[470]; 
    assign out[2599] = layer_0[4270] ^ layer_0[5023]; 
    assign out[2600] = ~layer_0[6275] | (layer_0[6275] & layer_0[7429]); 
    assign out[2601] = ~layer_0[5556] | (layer_0[5556] & layer_0[4543]); 
    assign out[2602] = layer_0[297]; 
    assign out[2603] = layer_0[7056]; 
    assign out[2604] = ~layer_0[4201]; 
    assign out[2605] = layer_0[2615] ^ layer_0[7654]; 
    assign out[2606] = layer_0[3585]; 
    assign out[2607] = ~(layer_0[2075] & layer_0[7925]); 
    assign out[2608] = ~(layer_0[4919] ^ layer_0[7870]); 
    assign out[2609] = layer_0[329] ^ layer_0[4403]; 
    assign out[2610] = ~layer_0[5176] | (layer_0[6467] & layer_0[5176]); 
    assign out[2611] = layer_0[544] & ~layer_0[414]; 
    assign out[2612] = ~(layer_0[3308] & layer_0[4563]); 
    assign out[2613] = layer_0[7713]; 
    assign out[2614] = ~(layer_0[6649] | layer_0[5647]); 
    assign out[2615] = ~(layer_0[1533] & layer_0[124]); 
    assign out[2616] = layer_0[36]; 
    assign out[2617] = ~layer_0[6412]; 
    assign out[2618] = layer_0[5642]; 
    assign out[2619] = layer_0[980] ^ layer_0[7602]; 
    assign out[2620] = ~layer_0[1307]; 
    assign out[2621] = layer_0[1875] ^ layer_0[2260]; 
    assign out[2622] = layer_0[6244]; 
    assign out[2623] = ~(layer_0[2173] | layer_0[3476]); 
    assign out[2624] = ~(layer_0[2414] & layer_0[660]); 
    assign out[2625] = ~(layer_0[718] & layer_0[650]); 
    assign out[2626] = ~layer_0[3275]; 
    assign out[2627] = ~(layer_0[299] ^ layer_0[1083]); 
    assign out[2628] = ~layer_0[4953] | (layer_0[4953] & layer_0[729]); 
    assign out[2629] = layer_0[1881] & layer_0[6217]; 
    assign out[2630] = ~(layer_0[6817] & layer_0[3504]); 
    assign out[2631] = ~layer_0[3820] | (layer_0[186] & layer_0[3820]); 
    assign out[2632] = layer_0[2301]; 
    assign out[2633] = layer_0[7838] ^ layer_0[2721]; 
    assign out[2634] = ~(layer_0[1784] ^ layer_0[1032]); 
    assign out[2635] = ~(layer_0[3898] & layer_0[1012]); 
    assign out[2636] = ~layer_0[3241] | (layer_0[5633] & layer_0[3241]); 
    assign out[2637] = layer_0[1402]; 
    assign out[2638] = ~(layer_0[6077] ^ layer_0[2859]); 
    assign out[2639] = layer_0[1585] | layer_0[6902]; 
    assign out[2640] = layer_0[6813] & ~layer_0[6697]; 
    assign out[2641] = layer_0[6599]; 
    assign out[2642] = layer_0[6820]; 
    assign out[2643] = ~layer_0[780]; 
    assign out[2644] = layer_0[6829]; 
    assign out[2645] = layer_0[2889]; 
    assign out[2646] = layer_0[2445]; 
    assign out[2647] = ~(layer_0[3282] & layer_0[5426]); 
    assign out[2648] = ~layer_0[7707] | (layer_0[7707] & layer_0[828]); 
    assign out[2649] = layer_0[2854] | layer_0[876]; 
    assign out[2650] = ~(layer_0[6057] ^ layer_0[6509]); 
    assign out[2651] = ~layer_0[5487]; 
    assign out[2652] = ~(layer_0[3999] ^ layer_0[3045]); 
    assign out[2653] = layer_0[7768] & ~layer_0[5540]; 
    assign out[2654] = ~(layer_0[7953] & layer_0[5331]); 
    assign out[2655] = ~layer_0[2813] | (layer_0[49] & layer_0[2813]); 
    assign out[2656] = ~(layer_0[4734] ^ layer_0[4044]); 
    assign out[2657] = layer_0[4170] & ~layer_0[1394]; 
    assign out[2658] = ~layer_0[6182] | (layer_0[6182] & layer_0[549]); 
    assign out[2659] = ~layer_0[345] | (layer_0[2910] & layer_0[345]); 
    assign out[2660] = ~(layer_0[2480] ^ layer_0[5566]); 
    assign out[2661] = ~layer_0[188]; 
    assign out[2662] = ~layer_0[6529] | (layer_0[7264] & layer_0[6529]); 
    assign out[2663] = layer_0[1670]; 
    assign out[2664] = ~(layer_0[1904] | layer_0[2826]); 
    assign out[2665] = ~layer_0[6539]; 
    assign out[2666] = ~layer_0[213]; 
    assign out[2667] = ~(layer_0[5237] ^ layer_0[803]); 
    assign out[2668] = layer_0[6292]; 
    assign out[2669] = layer_0[2573]; 
    assign out[2670] = ~layer_0[4466] | (layer_0[1337] & layer_0[4466]); 
    assign out[2671] = ~(layer_0[6849] & layer_0[3721]); 
    assign out[2672] = ~layer_0[5060] | (layer_0[5060] & layer_0[4050]); 
    assign out[2673] = ~(layer_0[654] & layer_0[6196]); 
    assign out[2674] = ~layer_0[3056]; 
    assign out[2675] = ~(layer_0[6898] & layer_0[3855]); 
    assign out[2676] = layer_0[538]; 
    assign out[2677] = ~layer_0[4640]; 
    assign out[2678] = ~layer_0[1478] | (layer_0[7618] & layer_0[1478]); 
    assign out[2679] = layer_0[1535] & ~layer_0[3180]; 
    assign out[2680] = ~layer_0[2842]; 
    assign out[2681] = layer_0[2049] ^ layer_0[5730]; 
    assign out[2682] = ~layer_0[612] | (layer_0[6763] & layer_0[612]); 
    assign out[2683] = ~layer_0[2145] | (layer_0[2145] & layer_0[2538]); 
    assign out[2684] = ~layer_0[5939]; 
    assign out[2685] = layer_0[5418] & ~layer_0[5921]; 
    assign out[2686] = layer_0[2780] & layer_0[4976]; 
    assign out[2687] = ~(layer_0[7400] ^ layer_0[931]); 
    assign out[2688] = ~layer_0[3933] | (layer_0[5747] & layer_0[3933]); 
    assign out[2689] = layer_0[1280]; 
    assign out[2690] = layer_0[3765]; 
    assign out[2691] = layer_0[5448] ^ layer_0[6852]; 
    assign out[2692] = layer_0[2293] ^ layer_0[3471]; 
    assign out[2693] = ~layer_0[5263]; 
    assign out[2694] = ~(layer_0[7597] ^ layer_0[1227]); 
    assign out[2695] = ~layer_0[863] | (layer_0[863] & layer_0[6519]); 
    assign out[2696] = ~layer_0[7037] | (layer_0[3420] & layer_0[7037]); 
    assign out[2697] = layer_0[1082] ^ layer_0[2254]; 
    assign out[2698] = ~layer_0[4691] | (layer_0[7734] & layer_0[4691]); 
    assign out[2699] = ~(layer_0[3322] & layer_0[6124]); 
    assign out[2700] = ~layer_0[1385]; 
    assign out[2701] = layer_0[5972]; 
    assign out[2702] = layer_0[1933]; 
    assign out[2703] = layer_0[3508]; 
    assign out[2704] = ~(layer_0[4132] ^ layer_0[5282]); 
    assign out[2705] = ~(layer_0[2164] & layer_0[2384]); 
    assign out[2706] = ~(layer_0[4288] ^ layer_0[6097]); 
    assign out[2707] = layer_0[4355]; 
    assign out[2708] = ~layer_0[1010]; 
    assign out[2709] = ~(layer_0[1891] ^ layer_0[6744]); 
    assign out[2710] = layer_0[7537] | layer_0[7373]; 
    assign out[2711] = ~layer_0[5737] | (layer_0[5737] & layer_0[3426]); 
    assign out[2712] = layer_0[6415]; 
    assign out[2713] = ~(layer_0[4231] ^ layer_0[7420]); 
    assign out[2714] = ~layer_0[4679] | (layer_0[4679] & layer_0[321]); 
    assign out[2715] = ~layer_0[7848] | (layer_0[2316] & layer_0[7848]); 
    assign out[2716] = layer_0[5920]; 
    assign out[2717] = ~(layer_0[7065] ^ layer_0[5066]); 
    assign out[2718] = layer_0[5689] ^ layer_0[39]; 
    assign out[2719] = ~layer_0[5044]; 
    assign out[2720] = ~layer_0[3698]; 
    assign out[2721] = ~(layer_0[1326] & layer_0[985]); 
    assign out[2722] = ~(layer_0[5502] & layer_0[4402]); 
    assign out[2723] = ~layer_0[6686] | (layer_0[6686] & layer_0[7797]); 
    assign out[2724] = ~(layer_0[4208] & layer_0[5777]); 
    assign out[2725] = ~(layer_0[6753] ^ layer_0[4122]); 
    assign out[2726] = ~layer_0[7685] | (layer_0[2499] & layer_0[7685]); 
    assign out[2727] = ~layer_0[7407] | (layer_0[7407] & layer_0[624]); 
    assign out[2728] = ~layer_0[2771]; 
    assign out[2729] = ~layer_0[6706]; 
    assign out[2730] = layer_0[3201]; 
    assign out[2731] = ~(layer_0[7183] & layer_0[177]); 
    assign out[2732] = layer_0[2748] ^ layer_0[7627]; 
    assign out[2733] = ~(layer_0[7443] & layer_0[719]); 
    assign out[2734] = layer_0[7697] | layer_0[1428]; 
    assign out[2735] = ~(layer_0[6578] ^ layer_0[2213]); 
    assign out[2736] = layer_0[2841]; 
    assign out[2737] = layer_0[4855] ^ layer_0[7334]; 
    assign out[2738] = ~layer_0[7232]; 
    assign out[2739] = ~(layer_0[5888] | layer_0[7540]); 
    assign out[2740] = layer_0[2271] ^ layer_0[6683]; 
    assign out[2741] = ~(layer_0[7635] & layer_0[7089]); 
    assign out[2742] = layer_0[4186] | layer_0[3938]; 
    assign out[2743] = ~(layer_0[1879] | layer_0[6898]); 
    assign out[2744] = ~(layer_0[685] ^ layer_0[4210]); 
    assign out[2745] = layer_0[2774] & layer_0[227]; 
    assign out[2746] = ~(layer_0[6504] | layer_0[7122]); 
    assign out[2747] = layer_0[7108] ^ layer_0[6466]; 
    assign out[2748] = ~layer_0[1823] | (layer_0[5153] & layer_0[1823]); 
    assign out[2749] = layer_0[2486] ^ layer_0[2477]; 
    assign out[2750] = ~layer_0[5321] | (layer_0[51] & layer_0[5321]); 
    assign out[2751] = ~(layer_0[3438] ^ layer_0[5086]); 
    assign out[2752] = ~(layer_0[3684] ^ layer_0[2953]); 
    assign out[2753] = ~layer_0[6109] | (layer_0[6109] & layer_0[1933]); 
    assign out[2754] = layer_0[2591] ^ layer_0[6993]; 
    assign out[2755] = layer_0[5600] & ~layer_0[6196]; 
    assign out[2756] = ~(layer_0[5969] ^ layer_0[5957]); 
    assign out[2757] = ~(layer_0[4958] ^ layer_0[1040]); 
    assign out[2758] = ~layer_0[1619]; 
    assign out[2759] = ~(layer_0[612] & layer_0[6523]); 
    assign out[2760] = ~layer_0[3094] | (layer_0[3094] & layer_0[897]); 
    assign out[2761] = ~layer_0[3733] | (layer_0[3733] & layer_0[2243]); 
    assign out[2762] = layer_0[3197] ^ layer_0[5686]; 
    assign out[2763] = ~layer_0[335]; 
    assign out[2764] = 1'b1; 
    assign out[2765] = layer_0[5938]; 
    assign out[2766] = ~layer_0[1828] | (layer_0[1828] & layer_0[840]); 
    assign out[2767] = ~layer_0[6327]; 
    assign out[2768] = ~layer_0[2901]; 
    assign out[2769] = ~layer_0[4486]; 
    assign out[2770] = layer_0[2717] ^ layer_0[6454]; 
    assign out[2771] = ~(layer_0[6534] ^ layer_0[526]); 
    assign out[2772] = ~layer_0[2959] | (layer_0[2959] & layer_0[6520]); 
    assign out[2773] = layer_0[6096]; 
    assign out[2774] = ~layer_0[261]; 
    assign out[2775] = ~(layer_0[7935] | layer_0[3710]); 
    assign out[2776] = ~layer_0[5879] | (layer_0[7073] & layer_0[5879]); 
    assign out[2777] = ~(layer_0[442] ^ layer_0[3688]); 
    assign out[2778] = ~(layer_0[594] ^ layer_0[4391]); 
    assign out[2779] = layer_0[425]; 
    assign out[2780] = ~layer_0[7908]; 
    assign out[2781] = layer_0[5701] ^ layer_0[487]; 
    assign out[2782] = layer_0[7929] | layer_0[5330]; 
    assign out[2783] = layer_0[6350] | layer_0[3873]; 
    assign out[2784] = ~layer_0[1926] | (layer_0[1926] & layer_0[1592]); 
    assign out[2785] = layer_0[5287] ^ layer_0[2387]; 
    assign out[2786] = ~(layer_0[1206] ^ layer_0[1408]); 
    assign out[2787] = ~(layer_0[613] & layer_0[6153]); 
    assign out[2788] = ~layer_0[4792]; 
    assign out[2789] = layer_0[3037] ^ layer_0[1698]; 
    assign out[2790] = layer_0[1540] ^ layer_0[2092]; 
    assign out[2791] = layer_0[7605] ^ layer_0[2448]; 
    assign out[2792] = ~layer_0[7098] | (layer_0[7098] & layer_0[7777]); 
    assign out[2793] = ~layer_0[7652]; 
    assign out[2794] = ~(layer_0[5018] ^ layer_0[101]); 
    assign out[2795] = layer_0[6839]; 
    assign out[2796] = ~(layer_0[7396] ^ layer_0[4866]); 
    assign out[2797] = layer_0[6730] | layer_0[5461]; 
    assign out[2798] = ~layer_0[1046]; 
    assign out[2799] = layer_0[4103]; 
    assign out[2800] = layer_0[3564] | layer_0[1242]; 
    assign out[2801] = ~layer_0[3632] | (layer_0[5793] & layer_0[3632]); 
    assign out[2802] = ~(layer_0[5539] ^ layer_0[7198]); 
    assign out[2803] = layer_0[6293] ^ layer_0[7503]; 
    assign out[2804] = ~layer_0[1177]; 
    assign out[2805] = layer_0[4064] ^ layer_0[5392]; 
    assign out[2806] = ~(layer_0[3987] ^ layer_0[3731]); 
    assign out[2807] = layer_0[1293] & layer_0[622]; 
    assign out[2808] = ~(layer_0[7436] & layer_0[781]); 
    assign out[2809] = ~layer_0[2373]; 
    assign out[2810] = layer_0[6622]; 
    assign out[2811] = ~(layer_0[4467] ^ layer_0[7430]); 
    assign out[2812] = ~layer_0[2905]; 
    assign out[2813] = layer_0[6068]; 
    assign out[2814] = layer_0[5121] & ~layer_0[19]; 
    assign out[2815] = ~layer_0[7076]; 
    assign out[2816] = ~(layer_0[1368] ^ layer_0[7124]); 
    assign out[2817] = layer_0[3424]; 
    assign out[2818] = layer_0[7981]; 
    assign out[2819] = ~layer_0[6125]; 
    assign out[2820] = layer_0[7710] & ~layer_0[6604]; 
    assign out[2821] = layer_0[4779]; 
    assign out[2822] = ~layer_0[2730] | (layer_0[1835] & layer_0[2730]); 
    assign out[2823] = ~(layer_0[5470] ^ layer_0[5108]); 
    assign out[2824] = ~layer_0[1313] | (layer_0[1116] & layer_0[1313]); 
    assign out[2825] = ~(layer_0[3616] ^ layer_0[7917]); 
    assign out[2826] = ~layer_0[1862] | (layer_0[1862] & layer_0[5623]); 
    assign out[2827] = layer_0[3160]; 
    assign out[2828] = ~layer_0[678]; 
    assign out[2829] = layer_0[1314]; 
    assign out[2830] = ~(layer_0[698] ^ layer_0[995]); 
    assign out[2831] = layer_0[5956] ^ layer_0[7409]; 
    assign out[2832] = ~(layer_0[7345] ^ layer_0[3178]); 
    assign out[2833] = ~(layer_0[7693] ^ layer_0[650]); 
    assign out[2834] = ~layer_0[419]; 
    assign out[2835] = ~(layer_0[7776] & layer_0[7573]); 
    assign out[2836] = layer_0[7601] ^ layer_0[6522]; 
    assign out[2837] = layer_0[3795] | layer_0[2745]; 
    assign out[2838] = ~(layer_0[86] & layer_0[1085]); 
    assign out[2839] = ~(layer_0[6270] ^ layer_0[3877]); 
    assign out[2840] = layer_0[6918]; 
    assign out[2841] = layer_0[2483] & layer_0[5488]; 
    assign out[2842] = ~layer_0[4146] | (layer_0[4146] & layer_0[3454]); 
    assign out[2843] = layer_0[3160] & ~layer_0[2828]; 
    assign out[2844] = ~(layer_0[6217] ^ layer_0[6772]); 
    assign out[2845] = ~(layer_0[7256] ^ layer_0[623]); 
    assign out[2846] = layer_0[2516] & ~layer_0[3169]; 
    assign out[2847] = ~(layer_0[7360] ^ layer_0[2371]); 
    assign out[2848] = ~layer_0[2914] | (layer_0[4811] & layer_0[2914]); 
    assign out[2849] = layer_0[1371] ^ layer_0[4046]; 
    assign out[2850] = ~layer_0[2893] | (layer_0[2893] & layer_0[4788]); 
    assign out[2851] = ~layer_0[2251] | (layer_0[2251] & layer_0[1302]); 
    assign out[2852] = ~layer_0[6115]; 
    assign out[2853] = layer_0[4502]; 
    assign out[2854] = ~(layer_0[7233] ^ layer_0[2855]); 
    assign out[2855] = layer_0[722] ^ layer_0[4352]; 
    assign out[2856] = ~(layer_0[7831] ^ layer_0[5909]); 
    assign out[2857] = ~layer_0[1504] | (layer_0[2368] & layer_0[1504]); 
    assign out[2858] = layer_0[1854] ^ layer_0[4754]; 
    assign out[2859] = layer_0[1766] & layer_0[4687]; 
    assign out[2860] = ~layer_0[5395] | (layer_0[5395] & layer_0[7136]); 
    assign out[2861] = layer_0[504] | layer_0[2802]; 
    assign out[2862] = ~layer_0[5548] | (layer_0[5548] & layer_0[2012]); 
    assign out[2863] = ~layer_0[536] | (layer_0[7032] & layer_0[536]); 
    assign out[2864] = ~layer_0[7342] | (layer_0[6012] & layer_0[7342]); 
    assign out[2865] = ~layer_0[4827]; 
    assign out[2866] = layer_0[2370] ^ layer_0[3993]; 
    assign out[2867] = layer_0[4304]; 
    assign out[2868] = layer_0[6424] | layer_0[7812]; 
    assign out[2869] = layer_0[2193] & ~layer_0[7051]; 
    assign out[2870] = layer_0[4285]; 
    assign out[2871] = layer_0[770]; 
    assign out[2872] = layer_0[6435] ^ layer_0[4762]; 
    assign out[2873] = ~(layer_0[2768] & layer_0[670]); 
    assign out[2874] = ~(layer_0[5698] ^ layer_0[4681]); 
    assign out[2875] = layer_0[6728] & layer_0[1293]; 
    assign out[2876] = ~(layer_0[1522] & layer_0[4598]); 
    assign out[2877] = ~(layer_0[2000] ^ layer_0[6654]); 
    assign out[2878] = ~(layer_0[4923] ^ layer_0[6897]); 
    assign out[2879] = layer_0[1975]; 
    assign out[2880] = layer_0[4279] & ~layer_0[1149]; 
    assign out[2881] = ~layer_0[301]; 
    assign out[2882] = layer_0[6538] ^ layer_0[3293]; 
    assign out[2883] = ~layer_0[7212] | (layer_0[4914] & layer_0[7212]); 
    assign out[2884] = layer_0[1019]; 
    assign out[2885] = layer_0[1881] & ~layer_0[7924]; 
    assign out[2886] = layer_0[2810]; 
    assign out[2887] = layer_0[3435] ^ layer_0[2471]; 
    assign out[2888] = layer_0[5967] ^ layer_0[54]; 
    assign out[2889] = ~layer_0[3709] | (layer_0[4101] & layer_0[3709]); 
    assign out[2890] = layer_0[6834] ^ layer_0[2930]; 
    assign out[2891] = ~(layer_0[3711] ^ layer_0[6229]); 
    assign out[2892] = layer_0[2956] ^ layer_0[5871]; 
    assign out[2893] = ~(layer_0[34] & layer_0[6498]); 
    assign out[2894] = layer_0[7346]; 
    assign out[2895] = ~(layer_0[4361] ^ layer_0[5708]); 
    assign out[2896] = layer_0[3353] ^ layer_0[2487]; 
    assign out[2897] = ~layer_0[472]; 
    assign out[2898] = ~(layer_0[2727] | layer_0[4724]); 
    assign out[2899] = ~(layer_0[1160] & layer_0[6708]); 
    assign out[2900] = ~layer_0[963] | (layer_0[527] & layer_0[963]); 
    assign out[2901] = layer_0[5483]; 
    assign out[2902] = ~layer_0[3912] | (layer_0[3912] & layer_0[1738]); 
    assign out[2903] = ~layer_0[5755] | (layer_0[5755] & layer_0[3366]); 
    assign out[2904] = layer_0[7181] ^ layer_0[351]; 
    assign out[2905] = ~layer_0[1732]; 
    assign out[2906] = ~layer_0[5596] | (layer_0[1929] & layer_0[5596]); 
    assign out[2907] = layer_0[5319] ^ layer_0[2454]; 
    assign out[2908] = ~(layer_0[2475] ^ layer_0[6804]); 
    assign out[2909] = ~layer_0[3675]; 
    assign out[2910] = ~layer_0[7918]; 
    assign out[2911] = layer_0[1186]; 
    assign out[2912] = ~layer_0[7224] | (layer_0[5662] & layer_0[7224]); 
    assign out[2913] = ~(layer_0[20] ^ layer_0[2896]); 
    assign out[2914] = layer_0[7011] ^ layer_0[6714]; 
    assign out[2915] = ~layer_0[2011] | (layer_0[2011] & layer_0[4255]); 
    assign out[2916] = ~layer_0[2940]; 
    assign out[2917] = layer_0[297]; 
    assign out[2918] = layer_0[3620] & ~layer_0[2284]; 
    assign out[2919] = layer_0[6845] | layer_0[1430]; 
    assign out[2920] = layer_0[493]; 
    assign out[2921] = layer_0[6907]; 
    assign out[2922] = layer_0[1202]; 
    assign out[2923] = layer_0[6381] ^ layer_0[4327]; 
    assign out[2924] = ~(layer_0[4878] | layer_0[1583]); 
    assign out[2925] = layer_0[112] ^ layer_0[7159]; 
    assign out[2926] = ~layer_0[4258] | (layer_0[6974] & layer_0[4258]); 
    assign out[2927] = ~layer_0[7803] | (layer_0[4193] & layer_0[7803]); 
    assign out[2928] = layer_0[4911] & ~layer_0[6382]; 
    assign out[2929] = ~(layer_0[6047] | layer_0[6869]); 
    assign out[2930] = ~(layer_0[3871] & layer_0[1495]); 
    assign out[2931] = ~layer_0[5745]; 
    assign out[2932] = ~(layer_0[7205] & layer_0[1142]); 
    assign out[2933] = layer_0[5156] ^ layer_0[2890]; 
    assign out[2934] = layer_0[4008]; 
    assign out[2935] = ~layer_0[6595] | (layer_0[6595] & layer_0[2511]); 
    assign out[2936] = layer_0[5677] ^ layer_0[6760]; 
    assign out[2937] = ~layer_0[7868] | (layer_0[7868] & layer_0[6998]); 
    assign out[2938] = ~layer_0[2168]; 
    assign out[2939] = ~(layer_0[2941] | layer_0[6100]); 
    assign out[2940] = ~layer_0[7276]; 
    assign out[2941] = ~(layer_0[4119] ^ layer_0[3949]); 
    assign out[2942] = layer_0[1043] ^ layer_0[5407]; 
    assign out[2943] = layer_0[5823] ^ layer_0[4618]; 
    assign out[2944] = ~layer_0[3092] | (layer_0[6953] & layer_0[3092]); 
    assign out[2945] = ~layer_0[4557]; 
    assign out[2946] = ~(layer_0[4061] ^ layer_0[2131]); 
    assign out[2947] = layer_0[3672]; 
    assign out[2948] = ~layer_0[6429] | (layer_0[479] & layer_0[6429]); 
    assign out[2949] = ~(layer_0[5771] ^ layer_0[4415]); 
    assign out[2950] = ~(layer_0[936] | layer_0[1321]); 
    assign out[2951] = layer_0[809]; 
    assign out[2952] = layer_0[3409]; 
    assign out[2953] = layer_0[2130] ^ layer_0[5666]; 
    assign out[2954] = ~layer_0[6371]; 
    assign out[2955] = ~layer_0[2801]; 
    assign out[2956] = layer_0[3381] ^ layer_0[5254]; 
    assign out[2957] = ~layer_0[2507]; 
    assign out[2958] = ~layer_0[4986]; 
    assign out[2959] = layer_0[1700]; 
    assign out[2960] = ~layer_0[7423] | (layer_0[7423] & layer_0[3678]); 
    assign out[2961] = ~(layer_0[1221] ^ layer_0[3450]); 
    assign out[2962] = ~layer_0[6302] | (layer_0[6302] & layer_0[6251]); 
    assign out[2963] = ~layer_0[5809] | (layer_0[5809] & layer_0[1052]); 
    assign out[2964] = layer_0[4153]; 
    assign out[2965] = ~layer_0[2468]; 
    assign out[2966] = ~layer_0[714] | (layer_0[714] & layer_0[7733]); 
    assign out[2967] = layer_0[4677]; 
    assign out[2968] = ~layer_0[1745]; 
    assign out[2969] = ~(layer_0[6723] & layer_0[593]); 
    assign out[2970] = layer_0[2388] ^ layer_0[1325]; 
    assign out[2971] = layer_0[2229] | layer_0[3797]; 
    assign out[2972] = layer_0[3614] | layer_0[3658]; 
    assign out[2973] = ~layer_0[4531]; 
    assign out[2974] = layer_0[7934] | layer_0[1284]; 
    assign out[2975] = layer_0[2309] ^ layer_0[2994]; 
    assign out[2976] = layer_0[473] | layer_0[7487]; 
    assign out[2977] = layer_0[5103] ^ layer_0[2034]; 
    assign out[2978] = layer_0[1270] ^ layer_0[37]; 
    assign out[2979] = layer_0[36] | layer_0[2194]; 
    assign out[2980] = layer_0[2991] | layer_0[1647]; 
    assign out[2981] = layer_0[2526]; 
    assign out[2982] = layer_0[7087] | layer_0[4537]; 
    assign out[2983] = ~layer_0[3719] | (layer_0[3719] & layer_0[6005]); 
    assign out[2984] = layer_0[416] & ~layer_0[207]; 
    assign out[2985] = layer_0[4586]; 
    assign out[2986] = layer_0[1059]; 
    assign out[2987] = layer_0[1710] ^ layer_0[4084]; 
    assign out[2988] = ~(layer_0[2756] ^ layer_0[2640]); 
    assign out[2989] = ~layer_0[7003] | (layer_0[7003] & layer_0[391]); 
    assign out[2990] = ~layer_0[7977] | (layer_0[1884] & layer_0[7977]); 
    assign out[2991] = layer_0[7103]; 
    assign out[2992] = layer_0[2844] | layer_0[7808]; 
    assign out[2993] = layer_0[1742] ^ layer_0[2437]; 
    assign out[2994] = layer_0[5813] & ~layer_0[4995]; 
    assign out[2995] = layer_0[1771]; 
    assign out[2996] = layer_0[5752] | layer_0[1079]; 
    assign out[2997] = layer_0[7781]; 
    assign out[2998] = ~(layer_0[614] & layer_0[5262]); 
    assign out[2999] = layer_0[5107] ^ layer_0[3885]; 
    assign out[3000] = layer_0[3761] | layer_0[3465]; 
    assign out[3001] = ~(layer_0[7678] | layer_0[5070]); 
    assign out[3002] = layer_0[7642] | layer_0[330]; 
    assign out[3003] = ~(layer_0[7391] ^ layer_0[6158]); 
    assign out[3004] = ~(layer_0[7559] & layer_0[6639]); 
    assign out[3005] = ~(layer_0[3349] ^ layer_0[6189]); 
    assign out[3006] = ~(layer_0[667] ^ layer_0[727]); 
    assign out[3007] = ~(layer_0[4615] ^ layer_0[5233]); 
    assign out[3008] = ~layer_0[1510] | (layer_0[4849] & layer_0[1510]); 
    assign out[3009] = ~(layer_0[6215] ^ layer_0[5749]); 
    assign out[3010] = layer_0[3326] ^ layer_0[829]; 
    assign out[3011] = ~(layer_0[2593] | layer_0[1119]); 
    assign out[3012] = ~layer_0[6551]; 
    assign out[3013] = ~(layer_0[4994] ^ layer_0[4577]); 
    assign out[3014] = ~layer_0[5607]; 
    assign out[3015] = ~layer_0[2073] | (layer_0[2073] & layer_0[4952]); 
    assign out[3016] = layer_0[3699] ^ layer_0[7795]; 
    assign out[3017] = layer_0[5186] | layer_0[254]; 
    assign out[3018] = layer_0[6149]; 
    assign out[3019] = layer_0[5279] | layer_0[4889]; 
    assign out[3020] = layer_0[7542] ^ layer_0[7425]; 
    assign out[3021] = ~layer_0[7453]; 
    assign out[3022] = ~layer_0[2264] | (layer_0[7992] & layer_0[2264]); 
    assign out[3023] = ~(layer_0[5131] ^ layer_0[113]); 
    assign out[3024] = ~layer_0[1343]; 
    assign out[3025] = ~(layer_0[1998] & layer_0[1589]); 
    assign out[3026] = ~layer_0[4088] | (layer_0[1824] & layer_0[4088]); 
    assign out[3027] = layer_0[6129] & ~layer_0[5881]; 
    assign out[3028] = layer_0[1323] ^ layer_0[7161]; 
    assign out[3029] = layer_0[7396] ^ layer_0[4005]; 
    assign out[3030] = layer_0[1040] ^ layer_0[5905]; 
    assign out[3031] = ~layer_0[3389] | (layer_0[3932] & layer_0[3389]); 
    assign out[3032] = ~(layer_0[275] ^ layer_0[1536]); 
    assign out[3033] = ~(layer_0[2833] ^ layer_0[4699]); 
    assign out[3034] = ~(layer_0[2578] & layer_0[3347]); 
    assign out[3035] = layer_0[850]; 
    assign out[3036] = ~(layer_0[5673] | layer_0[1898]); 
    assign out[3037] = layer_0[4134]; 
    assign out[3038] = ~(layer_0[5901] | layer_0[1734]); 
    assign out[3039] = ~layer_0[368]; 
    assign out[3040] = layer_0[3044] ^ layer_0[417]; 
    assign out[3041] = ~layer_0[1292] | (layer_0[5161] & layer_0[1292]); 
    assign out[3042] = layer_0[575] ^ layer_0[7492]; 
    assign out[3043] = ~layer_0[2782]; 
    assign out[3044] = layer_0[3381] ^ layer_0[3028]; 
    assign out[3045] = ~(layer_0[1970] | layer_0[5035]); 
    assign out[3046] = ~layer_0[737] | (layer_0[85] & layer_0[737]); 
    assign out[3047] = ~layer_0[489]; 
    assign out[3048] = ~layer_0[533]; 
    assign out[3049] = ~layer_0[7681]; 
    assign out[3050] = ~layer_0[7914]; 
    assign out[3051] = ~(layer_0[5310] | layer_0[5811]); 
    assign out[3052] = ~layer_0[1882] | (layer_0[1882] & layer_0[3880]); 
    assign out[3053] = layer_0[456] | layer_0[4690]; 
    assign out[3054] = ~layer_0[4425]; 
    assign out[3055] = layer_0[7157] & ~layer_0[6436]; 
    assign out[3056] = ~(layer_0[6399] ^ layer_0[3976]); 
    assign out[3057] = layer_0[5075] | layer_0[862]; 
    assign out[3058] = layer_0[2070]; 
    assign out[3059] = ~layer_0[1571] | (layer_0[1571] & layer_0[1454]); 
    assign out[3060] = layer_0[607]; 
    assign out[3061] = ~(layer_0[5638] ^ layer_0[5357]); 
    assign out[3062] = ~layer_0[5159]; 
    assign out[3063] = ~(layer_0[818] ^ layer_0[4164]); 
    assign out[3064] = ~layer_0[2832]; 
    assign out[3065] = ~layer_0[2331]; 
    assign out[3066] = ~(layer_0[1059] | layer_0[1279]); 
    assign out[3067] = layer_0[423] ^ layer_0[2474]; 
    assign out[3068] = ~(layer_0[7883] ^ layer_0[851]); 
    assign out[3069] = ~(layer_0[5599] & layer_0[60]); 
    assign out[3070] = layer_0[3280] ^ layer_0[312]; 
    assign out[3071] = ~layer_0[7807]; 
    assign out[3072] = layer_0[7861] ^ layer_0[7580]; 
    assign out[3073] = ~layer_0[3645] | (layer_0[3645] & layer_0[3556]); 
    assign out[3074] = ~(layer_0[7420] ^ layer_0[3250]); 
    assign out[3075] = layer_0[6260] & ~layer_0[2384]; 
    assign out[3076] = ~layer_0[3474]; 
    assign out[3077] = ~(layer_0[5692] & layer_0[5241]); 
    assign out[3078] = layer_0[1919] ^ layer_0[2265]; 
    assign out[3079] = layer_0[2392] ^ layer_0[3581]; 
    assign out[3080] = ~layer_0[627] | (layer_0[627] & layer_0[2605]); 
    assign out[3081] = layer_0[1656] ^ layer_0[3808]; 
    assign out[3082] = layer_0[5733] ^ layer_0[6506]; 
    assign out[3083] = layer_0[6735]; 
    assign out[3084] = ~(layer_0[5490] ^ layer_0[7850]); 
    assign out[3085] = ~(layer_0[4416] ^ layer_0[7758]); 
    assign out[3086] = layer_0[2775] & layer_0[3092]; 
    assign out[3087] = ~(layer_0[6773] ^ layer_0[1980]); 
    assign out[3088] = ~layer_0[7990]; 
    assign out[3089] = layer_0[7160] | layer_0[1703]; 
    assign out[3090] = ~(layer_0[1782] ^ layer_0[201]); 
    assign out[3091] = ~(layer_0[6532] ^ layer_0[6035]); 
    assign out[3092] = ~(layer_0[7796] ^ layer_0[7901]); 
    assign out[3093] = ~(layer_0[6192] | layer_0[1025]); 
    assign out[3094] = ~layer_0[1856]; 
    assign out[3095] = layer_0[5215] ^ layer_0[7191]; 
    assign out[3096] = layer_0[6782]; 
    assign out[3097] = ~(layer_0[6016] ^ layer_0[4517]); 
    assign out[3098] = layer_0[2062]; 
    assign out[3099] = ~layer_0[4941] | (layer_0[4941] & layer_0[6050]); 
    assign out[3100] = ~layer_0[3320] | (layer_0[3055] & layer_0[3320]); 
    assign out[3101] = ~(layer_0[983] & layer_0[4421]); 
    assign out[3102] = ~(layer_0[1381] ^ layer_0[3082]); 
    assign out[3103] = ~(layer_0[6203] ^ layer_0[2128]); 
    assign out[3104] = layer_0[7226] | layer_0[543]; 
    assign out[3105] = ~(layer_0[1792] ^ layer_0[133]); 
    assign out[3106] = ~layer_0[4213]; 
    assign out[3107] = layer_0[5966]; 
    assign out[3108] = ~(layer_0[7384] ^ layer_0[4014]); 
    assign out[3109] = layer_0[104]; 
    assign out[3110] = layer_0[1984] & ~layer_0[2936]; 
    assign out[3111] = layer_0[5381] | layer_0[1432]; 
    assign out[3112] = ~(layer_0[3509] ^ layer_0[4581]); 
    assign out[3113] = layer_0[2508] ^ layer_0[2038]; 
    assign out[3114] = ~layer_0[4117] | (layer_0[2617] & layer_0[4117]); 
    assign out[3115] = ~layer_0[3196]; 
    assign out[3116] = layer_0[4242] ^ layer_0[2843]; 
    assign out[3117] = layer_0[97] | layer_0[4993]; 
    assign out[3118] = layer_0[2008] ^ layer_0[3017]; 
    assign out[3119] = ~(layer_0[6127] | layer_0[3742]); 
    assign out[3120] = ~(layer_0[4751] ^ layer_0[1392]); 
    assign out[3121] = layer_0[4471] & ~layer_0[527]; 
    assign out[3122] = layer_0[2966]; 
    assign out[3123] = ~(layer_0[2857] ^ layer_0[2447]); 
    assign out[3124] = layer_0[6209] & layer_0[5397]; 
    assign out[3125] = layer_0[6225] ^ layer_0[3735]; 
    assign out[3126] = ~(layer_0[1867] ^ layer_0[4494]); 
    assign out[3127] = ~(layer_0[3795] ^ layer_0[5008]); 
    assign out[3128] = ~(layer_0[6265] ^ layer_0[1650]); 
    assign out[3129] = layer_0[3827] ^ layer_0[414]; 
    assign out[3130] = ~(layer_0[6592] & layer_0[7969]); 
    assign out[3131] = layer_0[3851] ^ layer_0[6656]; 
    assign out[3132] = ~(layer_0[7379] | layer_0[4805]); 
    assign out[3133] = layer_0[7835] ^ layer_0[4756]; 
    assign out[3134] = layer_0[4799] ^ layer_0[4315]; 
    assign out[3135] = layer_0[3299] & ~layer_0[5316]; 
    assign out[3136] = layer_0[3225] ^ layer_0[6237]; 
    assign out[3137] = layer_0[4723]; 
    assign out[3138] = ~(layer_0[6156] ^ layer_0[4012]); 
    assign out[3139] = ~(layer_0[1519] | layer_0[153]); 
    assign out[3140] = layer_0[5958]; 
    assign out[3141] = layer_0[587]; 
    assign out[3142] = ~(layer_0[191] & layer_0[187]); 
    assign out[3143] = layer_0[3210] & layer_0[3590]; 
    assign out[3144] = ~layer_0[7476]; 
    assign out[3145] = layer_0[7593] ^ layer_0[6603]; 
    assign out[3146] = layer_0[1124] ^ layer_0[349]; 
    assign out[3147] = layer_0[273] & ~layer_0[5009]; 
    assign out[3148] = layer_0[4109]; 
    assign out[3149] = layer_0[7508] ^ layer_0[205]; 
    assign out[3150] = layer_0[6101] & ~layer_0[5781]; 
    assign out[3151] = layer_0[5958] & layer_0[528]; 
    assign out[3152] = ~(layer_0[6209] ^ layer_0[3395]); 
    assign out[3153] = ~(layer_0[6688] ^ layer_0[4459]); 
    assign out[3154] = layer_0[424] & ~layer_0[6848]; 
    assign out[3155] = ~(layer_0[6262] & layer_0[1080]); 
    assign out[3156] = ~layer_0[4404]; 
    assign out[3157] = ~layer_0[2726] | (layer_0[2726] & layer_0[925]); 
    assign out[3158] = layer_0[6673]; 
    assign out[3159] = layer_0[6239] | layer_0[2094]; 
    assign out[3160] = layer_0[3022] ^ layer_0[2463]; 
    assign out[3161] = layer_0[982] ^ layer_0[2256]; 
    assign out[3162] = ~(layer_0[6715] ^ layer_0[1316]); 
    assign out[3163] = layer_0[3256] | layer_0[1511]; 
    assign out[3164] = layer_0[2067] ^ layer_0[4501]; 
    assign out[3165] = ~(layer_0[7705] ^ layer_0[6151]); 
    assign out[3166] = layer_0[3229]; 
    assign out[3167] = ~layer_0[2241] | (layer_0[2241] & layer_0[4206]); 
    assign out[3168] = ~(layer_0[1377] ^ layer_0[2212]); 
    assign out[3169] = layer_0[6114] ^ layer_0[6284]; 
    assign out[3170] = ~(layer_0[6411] ^ layer_0[5661]); 
    assign out[3171] = layer_0[1214]; 
    assign out[3172] = layer_0[6116] & ~layer_0[1889]; 
    assign out[3173] = layer_0[3861] | layer_0[1509]; 
    assign out[3174] = layer_0[4268] & ~layer_0[5786]; 
    assign out[3175] = ~(layer_0[7671] ^ layer_0[1097]); 
    assign out[3176] = ~(layer_0[576] ^ layer_0[2492]); 
    assign out[3177] = layer_0[4801]; 
    assign out[3178] = ~(layer_0[6816] ^ layer_0[5497]); 
    assign out[3179] = layer_0[1872] ^ layer_0[2141]; 
    assign out[3180] = layer_0[4524] ^ layer_0[1467]; 
    assign out[3181] = ~(layer_0[452] ^ layer_0[5825]); 
    assign out[3182] = layer_0[7209] & layer_0[5448]; 
    assign out[3183] = ~(layer_0[2013] | layer_0[3948]); 
    assign out[3184] = ~(layer_0[4674] ^ layer_0[6620]); 
    assign out[3185] = ~(layer_0[3155] ^ layer_0[115]); 
    assign out[3186] = ~(layer_0[2087] ^ layer_0[4513]); 
    assign out[3187] = ~(layer_0[135] ^ layer_0[1688]); 
    assign out[3188] = ~(layer_0[254] ^ layer_0[2055]); 
    assign out[3189] = ~layer_0[6470] | (layer_0[3205] & layer_0[6470]); 
    assign out[3190] = layer_0[7104] ^ layer_0[1028]; 
    assign out[3191] = layer_0[7828] & ~layer_0[3891]; 
    assign out[3192] = ~layer_0[4896] | (layer_0[127] & layer_0[4896]); 
    assign out[3193] = ~layer_0[3466]; 
    assign out[3194] = layer_0[7305] & ~layer_0[3207]; 
    assign out[3195] = layer_0[2219]; 
    assign out[3196] = ~layer_0[1978] | (layer_0[5518] & layer_0[1978]); 
    assign out[3197] = ~(layer_0[6889] ^ layer_0[327]); 
    assign out[3198] = layer_0[3460] ^ layer_0[3043]; 
    assign out[3199] = layer_0[5284] ^ layer_0[2131]; 
    assign out[3200] = ~layer_0[6655] | (layer_0[1426] & layer_0[6655]); 
    assign out[3201] = ~(layer_0[7404] & layer_0[2277]); 
    assign out[3202] = ~(layer_0[5347] | layer_0[6876]); 
    assign out[3203] = layer_0[1762]; 
    assign out[3204] = layer_0[3562] ^ layer_0[1571]; 
    assign out[3205] = layer_0[7309]; 
    assign out[3206] = ~layer_0[5225] | (layer_0[2912] & layer_0[5225]); 
    assign out[3207] = layer_0[1851] | layer_0[5680]; 
    assign out[3208] = layer_0[6792] & ~layer_0[7335]; 
    assign out[3209] = ~(layer_0[3624] ^ layer_0[4374]); 
    assign out[3210] = ~(layer_0[2672] & layer_0[5364]); 
    assign out[3211] = layer_0[3754]; 
    assign out[3212] = ~(layer_0[1216] ^ layer_0[5920]); 
    assign out[3213] = ~(layer_0[5423] ^ layer_0[1833]); 
    assign out[3214] = layer_0[6640] ^ layer_0[930]; 
    assign out[3215] = layer_0[6566] ^ layer_0[4442]; 
    assign out[3216] = layer_0[5550] | layer_0[2971]; 
    assign out[3217] = ~layer_0[5050] | (layer_0[5050] & layer_0[3111]); 
    assign out[3218] = layer_0[7872] ^ layer_0[6569]; 
    assign out[3219] = ~(layer_0[1481] ^ layer_0[2253]); 
    assign out[3220] = ~(layer_0[4600] | layer_0[3343]); 
    assign out[3221] = ~layer_0[3360] | (layer_0[3360] & layer_0[6914]); 
    assign out[3222] = ~(layer_0[1027] & layer_0[4565]); 
    assign out[3223] = layer_0[3559] & layer_0[528]; 
    assign out[3224] = layer_0[7898] ^ layer_0[6722]; 
    assign out[3225] = ~(layer_0[6878] ^ layer_0[1406]); 
    assign out[3226] = layer_0[1338]; 
    assign out[3227] = layer_0[4607] ^ layer_0[4636]; 
    assign out[3228] = ~layer_0[5528] | (layer_0[2028] & layer_0[5528]); 
    assign out[3229] = ~layer_0[5986]; 
    assign out[3230] = ~layer_0[7744] | (layer_0[7744] & layer_0[6306]); 
    assign out[3231] = ~(layer_0[4408] ^ layer_0[1135]); 
    assign out[3232] = layer_0[7888] ^ layer_0[1155]; 
    assign out[3233] = ~(layer_0[4893] ^ layer_0[5951]); 
    assign out[3234] = ~(layer_0[3182] ^ layer_0[1913]); 
    assign out[3235] = layer_0[161] ^ layer_0[4868]; 
    assign out[3236] = ~layer_0[5179] | (layer_0[5179] & layer_0[2635]); 
    assign out[3237] = layer_0[6448] & ~layer_0[6540]; 
    assign out[3238] = ~(layer_0[1549] ^ layer_0[4497]); 
    assign out[3239] = ~(layer_0[6265] ^ layer_0[3895]); 
    assign out[3240] = layer_0[174] ^ layer_0[5047]; 
    assign out[3241] = layer_0[2433] ^ layer_0[205]; 
    assign out[3242] = layer_0[2348] | layer_0[177]; 
    assign out[3243] = layer_0[6905] ^ layer_0[4939]; 
    assign out[3244] = layer_0[454] ^ layer_0[5048]; 
    assign out[3245] = ~(layer_0[6966] ^ layer_0[6628]); 
    assign out[3246] = ~layer_0[2641] | (layer_0[2641] & layer_0[5903]); 
    assign out[3247] = ~(layer_0[2444] ^ layer_0[196]); 
    assign out[3248] = layer_0[1902] ^ layer_0[2332]; 
    assign out[3249] = ~(layer_0[2502] & layer_0[2047]); 
    assign out[3250] = layer_0[2972] ^ layer_0[3038]; 
    assign out[3251] = ~(layer_0[2479] ^ layer_0[6330]); 
    assign out[3252] = layer_0[3775] & ~layer_0[6993]; 
    assign out[3253] = ~layer_0[2950] | (layer_0[2950] & layer_0[3911]); 
    assign out[3254] = ~(layer_0[4406] ^ layer_0[6274]); 
    assign out[3255] = ~(layer_0[728] ^ layer_0[1458]); 
    assign out[3256] = ~layer_0[204]; 
    assign out[3257] = layer_0[5484]; 
    assign out[3258] = layer_0[6941] ^ layer_0[2103]; 
    assign out[3259] = ~(layer_0[7199] & layer_0[7548]); 
    assign out[3260] = layer_0[7258] & layer_0[1658]; 
    assign out[3261] = layer_0[7172] ^ layer_0[4514]; 
    assign out[3262] = ~(layer_0[7570] ^ layer_0[5906]); 
    assign out[3263] = ~(layer_0[260] & layer_0[2418]); 
    assign out[3264] = ~layer_0[1665]; 
    assign out[3265] = layer_0[1934] ^ layer_0[1918]; 
    assign out[3266] = layer_0[2659] ^ layer_0[7364]; 
    assign out[3267] = layer_0[3561] ^ layer_0[5640]; 
    assign out[3268] = ~(layer_0[5898] ^ layer_0[5197]); 
    assign out[3269] = layer_0[4624] ^ layer_0[706]; 
    assign out[3270] = layer_0[6597] & ~layer_0[2604]; 
    assign out[3271] = ~(layer_0[6620] ^ layer_0[1656]); 
    assign out[3272] = ~(layer_0[2037] ^ layer_0[4891]); 
    assign out[3273] = ~layer_0[3770] | (layer_0[1150] & layer_0[3770]); 
    assign out[3274] = ~layer_0[5982]; 
    assign out[3275] = ~layer_0[2112] | (layer_0[2112] & layer_0[7646]); 
    assign out[3276] = layer_0[5352] & layer_0[4170]; 
    assign out[3277] = ~(layer_0[5042] ^ layer_0[5743]); 
    assign out[3278] = ~(layer_0[1089] ^ layer_0[3631]); 
    assign out[3279] = layer_0[7621] & ~layer_0[3700]; 
    assign out[3280] = layer_0[576] ^ layer_0[6021]; 
    assign out[3281] = layer_0[5027] ^ layer_0[233]; 
    assign out[3282] = ~layer_0[6212] | (layer_0[4512] & layer_0[6212]); 
    assign out[3283] = layer_0[3199]; 
    assign out[3284] = ~(layer_0[402] ^ layer_0[766]); 
    assign out[3285] = layer_0[5298] ^ layer_0[3076]; 
    assign out[3286] = ~(layer_0[7684] ^ layer_0[7886]); 
    assign out[3287] = ~(layer_0[1471] ^ layer_0[7241]); 
    assign out[3288] = layer_0[7817] ^ layer_0[4179]; 
    assign out[3289] = layer_0[2700]; 
    assign out[3290] = ~(layer_0[3212] ^ layer_0[5704]); 
    assign out[3291] = layer_0[3534] ^ layer_0[7979]; 
    assign out[3292] = ~layer_0[6250] | (layer_0[6250] & layer_0[2439]); 
    assign out[3293] = layer_0[1062] | layer_0[7135]; 
    assign out[3294] = ~layer_0[7824] | (layer_0[7824] & layer_0[6395]); 
    assign out[3295] = ~layer_0[6720]; 
    assign out[3296] = layer_0[7485] ^ layer_0[6996]; 
    assign out[3297] = layer_0[1497]; 
    assign out[3298] = ~(layer_0[6528] & layer_0[7483]); 
    assign out[3299] = layer_0[6526] ^ layer_0[7023]; 
    assign out[3300] = ~(layer_0[2687] ^ layer_0[1569]); 
    assign out[3301] = ~(layer_0[6483] ^ layer_0[3968]); 
    assign out[3302] = layer_0[4967] ^ layer_0[6252]; 
    assign out[3303] = ~(layer_0[2246] & layer_0[2378]); 
    assign out[3304] = layer_0[2334] ^ layer_0[6019]; 
    assign out[3305] = ~(layer_0[4919] ^ layer_0[484]); 
    assign out[3306] = layer_0[3049]; 
    assign out[3307] = ~(layer_0[5360] ^ layer_0[3735]); 
    assign out[3308] = ~layer_0[1156] | (layer_0[1156] & layer_0[6161]); 
    assign out[3309] = layer_0[1246] ^ layer_0[2940]; 
    assign out[3310] = layer_0[919] ^ layer_0[6864]; 
    assign out[3311] = layer_0[2159]; 
    assign out[3312] = layer_0[6786]; 
    assign out[3313] = ~(layer_0[7788] ^ layer_0[4920]); 
    assign out[3314] = ~(layer_0[5090] ^ layer_0[4948]); 
    assign out[3315] = ~(layer_0[1281] ^ layer_0[2156]); 
    assign out[3316] = layer_0[3] | layer_0[3511]; 
    assign out[3317] = layer_0[3392]; 
    assign out[3318] = layer_0[1095] ^ layer_0[6073]; 
    assign out[3319] = ~(layer_0[61] ^ layer_0[3024]); 
    assign out[3320] = layer_0[3432] ^ layer_0[6818]; 
    assign out[3321] = layer_0[2251]; 
    assign out[3322] = layer_0[5842] ^ layer_0[423]; 
    assign out[3323] = ~layer_0[4905] | (layer_0[216] & layer_0[4905]); 
    assign out[3324] = layer_0[1637] ^ layer_0[84]; 
    assign out[3325] = layer_0[7288] ^ layer_0[4774]; 
    assign out[3326] = ~(layer_0[6437] ^ layer_0[6432]); 
    assign out[3327] = ~layer_0[3067]; 
    assign out[3328] = 1'b1; 
    assign out[3329] = layer_0[7014] ^ layer_0[2767]; 
    assign out[3330] = ~layer_0[3304]; 
    assign out[3331] = layer_0[209]; 
    assign out[3332] = layer_0[6222] ^ layer_0[7823]; 
    assign out[3333] = ~(layer_0[7246] & layer_0[6029]); 
    assign out[3334] = layer_0[3244] & ~layer_0[4491]; 
    assign out[3335] = ~layer_0[4611]; 
    assign out[3336] = layer_0[2777] ^ layer_0[1892]; 
    assign out[3337] = layer_0[6071] | layer_0[5597]; 
    assign out[3338] = ~(layer_0[3003] ^ layer_0[1617]); 
    assign out[3339] = ~(layer_0[2662] ^ layer_0[373]); 
    assign out[3340] = layer_0[2590] ^ layer_0[7012]; 
    assign out[3341] = ~(layer_0[7973] ^ layer_0[2421]); 
    assign out[3342] = ~(layer_0[4019] & layer_0[2315]); 
    assign out[3343] = layer_0[2299] ^ layer_0[3115]; 
    assign out[3344] = ~(layer_0[1157] ^ layer_0[2350]); 
    assign out[3345] = layer_0[117]; 
    assign out[3346] = layer_0[3149] & layer_0[1154]; 
    assign out[3347] = ~layer_0[7610]; 
    assign out[3348] = layer_0[434] ^ layer_0[170]; 
    assign out[3349] = layer_0[3242] | layer_0[6477]; 
    assign out[3350] = ~(layer_0[3104] ^ layer_0[465]); 
    assign out[3351] = ~(layer_0[4841] | layer_0[483]); 
    assign out[3352] = ~(layer_0[682] ^ layer_0[1649]); 
    assign out[3353] = ~layer_0[280]; 
    assign out[3354] = ~layer_0[3802] | (layer_0[3802] & layer_0[1350]); 
    assign out[3355] = ~(layer_0[41] | layer_0[2580]); 
    assign out[3356] = ~(layer_0[3341] ^ layer_0[7608]); 
    assign out[3357] = layer_0[646] & ~layer_0[1812]; 
    assign out[3358] = ~layer_0[3714] | (layer_0[3714] & layer_0[4619]); 
    assign out[3359] = ~layer_0[98]; 
    assign out[3360] = layer_0[325] ^ layer_0[1989]; 
    assign out[3361] = layer_0[6499] ^ layer_0[1100]; 
    assign out[3362] = ~(layer_0[630] ^ layer_0[160]); 
    assign out[3363] = layer_0[472] ^ layer_0[6090]; 
    assign out[3364] = ~(layer_0[6444] ^ layer_0[4861]); 
    assign out[3365] = ~layer_0[5778] | (layer_0[5778] & layer_0[1823]); 
    assign out[3366] = ~(layer_0[6870] ^ layer_0[7447]); 
    assign out[3367] = ~(layer_0[1712] ^ layer_0[325]); 
    assign out[3368] = ~layer_0[3097]; 
    assign out[3369] = ~(layer_0[1023] ^ layer_0[7876]); 
    assign out[3370] = layer_0[3768] ^ layer_0[4885]; 
    assign out[3371] = ~(layer_0[193] & layer_0[3472]); 
    assign out[3372] = ~(layer_0[4135] ^ layer_0[5310]); 
    assign out[3373] = layer_0[2171] ^ layer_0[7072]; 
    assign out[3374] = ~(layer_0[6616] ^ layer_0[4847]); 
    assign out[3375] = layer_0[901] ^ layer_0[7704]; 
    assign out[3376] = layer_0[5204]; 
    assign out[3377] = layer_0[4968] ^ layer_0[304]; 
    assign out[3378] = ~(layer_0[5127] & layer_0[7045]); 
    assign out[3379] = ~layer_0[3131]; 
    assign out[3380] = layer_0[7488] & ~layer_0[6374]; 
    assign out[3381] = layer_0[5592] ^ layer_0[2503]; 
    assign out[3382] = ~layer_0[2121] | (layer_0[2121] & layer_0[3660]); 
    assign out[3383] = layer_0[5261] ^ layer_0[939]; 
    assign out[3384] = ~layer_0[4369] | (layer_0[147] & layer_0[4369]); 
    assign out[3385] = layer_0[2275] ^ layer_0[1465]; 
    assign out[3386] = layer_0[2467]; 
    assign out[3387] = ~(layer_0[1396] ^ layer_0[2051]); 
    assign out[3388] = layer_0[3995] ^ layer_0[7125]; 
    assign out[3389] = layer_0[3218] ^ layer_0[3007]; 
    assign out[3390] = ~(layer_0[581] ^ layer_0[5286]); 
    assign out[3391] = ~(layer_0[2216] & layer_0[3557]); 
    assign out[3392] = layer_0[7154] & layer_0[880]; 
    assign out[3393] = ~(layer_0[2554] ^ layer_0[5754]); 
    assign out[3394] = layer_0[6249]; 
    assign out[3395] = layer_0[1106] ^ layer_0[992]; 
    assign out[3396] = layer_0[4510] | layer_0[4967]; 
    assign out[3397] = layer_0[7911] ^ layer_0[3333]; 
    assign out[3398] = layer_0[3365] ^ layer_0[4633]; 
    assign out[3399] = layer_0[5721]; 
    assign out[3400] = ~(layer_0[4487] | layer_0[1651]); 
    assign out[3401] = layer_0[7348] & ~layer_0[1410]; 
    assign out[3402] = layer_0[6912]; 
    assign out[3403] = ~(layer_0[7363] ^ layer_0[6712]); 
    assign out[3404] = layer_0[4354]; 
    assign out[3405] = layer_0[762]; 
    assign out[3406] = ~layer_0[2995] | (layer_0[3544] & layer_0[2995]); 
    assign out[3407] = layer_0[5978] ^ layer_0[5545]; 
    assign out[3408] = layer_0[4798] & ~layer_0[6596]; 
    assign out[3409] = ~layer_0[2706]; 
    assign out[3410] = layer_0[2628] ^ layer_0[1225]; 
    assign out[3411] = layer_0[3799] | layer_0[2957]; 
    assign out[3412] = layer_0[5643] ^ layer_0[3933]; 
    assign out[3413] = layer_0[7892] ^ layer_0[7193]; 
    assign out[3414] = ~(layer_0[4721] | layer_0[1473]); 
    assign out[3415] = layer_0[5240] & ~layer_0[6772]; 
    assign out[3416] = layer_0[409] ^ layer_0[4562]; 
    assign out[3417] = layer_0[5045] & ~layer_0[1902]; 
    assign out[3418] = ~layer_0[1635]; 
    assign out[3419] = ~layer_0[4388]; 
    assign out[3420] = ~layer_0[1364] | (layer_0[1364] & layer_0[5621]); 
    assign out[3421] = ~layer_0[6892] | (layer_0[2884] & layer_0[6892]); 
    assign out[3422] = ~(layer_0[7664] ^ layer_0[5725]); 
    assign out[3423] = ~(layer_0[1667] ^ layer_0[2804]); 
    assign out[3424] = layer_0[5918] ^ layer_0[2457]; 
    assign out[3425] = 1'b1; 
    assign out[3426] = layer_0[1260] ^ layer_0[1976]; 
    assign out[3427] = ~(layer_0[3479] & layer_0[5537]); 
    assign out[3428] = layer_0[4180] ^ layer_0[396]; 
    assign out[3429] = ~(layer_0[4924] ^ layer_0[4065]); 
    assign out[3430] = layer_0[1000] ^ layer_0[5439]; 
    assign out[3431] = ~layer_0[7606]; 
    assign out[3432] = ~layer_0[1640] | (layer_0[1240] & layer_0[1640]); 
    assign out[3433] = layer_0[2690] ^ layer_0[1296]; 
    assign out[3434] = ~(layer_0[7477] ^ layer_0[5433]); 
    assign out[3435] = ~(layer_0[2438] ^ layer_0[1545]); 
    assign out[3436] = ~(layer_0[5326] ^ layer_0[655]); 
    assign out[3437] = layer_0[7170] & ~layer_0[6911]; 
    assign out[3438] = ~(layer_0[3479] ^ layer_0[445]); 
    assign out[3439] = ~(layer_0[5659] ^ layer_0[3706]); 
    assign out[3440] = layer_0[4159] & layer_0[2786]; 
    assign out[3441] = layer_0[448] | layer_0[2405]; 
    assign out[3442] = layer_0[3446] ^ layer_0[6609]; 
    assign out[3443] = ~(layer_0[1579] ^ layer_0[6566]); 
    assign out[3444] = ~layer_0[1860]; 
    assign out[3445] = layer_0[4262] ^ layer_0[5807]; 
    assign out[3446] = layer_0[2260] ^ layer_0[7569]; 
    assign out[3447] = layer_0[7840] | layer_0[5456]; 
    assign out[3448] = ~(layer_0[310] & layer_0[5231]); 
    assign out[3449] = ~layer_0[1283]; 
    assign out[3450] = ~layer_0[284] | (layer_0[284] & layer_0[2001]); 
    assign out[3451] = ~(layer_0[4001] ^ layer_0[4320]); 
    assign out[3452] = layer_0[1175]; 
    assign out[3453] = ~layer_0[1344]; 
    assign out[3454] = layer_0[1793]; 
    assign out[3455] = ~(layer_0[474] ^ layer_0[7294]); 
    assign out[3456] = ~layer_0[3667] | (layer_0[3667] & layer_0[605]); 
    assign out[3457] = layer_0[6213] ^ layer_0[4246]; 
    assign out[3458] = ~(layer_0[486] ^ layer_0[4859]); 
    assign out[3459] = layer_0[2716] | layer_0[3812]; 
    assign out[3460] = ~layer_0[3072] | (layer_0[4493] & layer_0[3072]); 
    assign out[3461] = layer_0[7842]; 
    assign out[3462] = ~(layer_0[28] ^ layer_0[4711]); 
    assign out[3463] = layer_0[6207] & layer_0[6497]; 
    assign out[3464] = ~(layer_0[3412] ^ layer_0[4737]); 
    assign out[3465] = ~layer_0[4554] | (layer_0[5338] & layer_0[4554]); 
    assign out[3466] = ~layer_0[6061] | (layer_0[3680] & layer_0[6061]); 
    assign out[3467] = layer_0[4909] ^ layer_0[3290]; 
    assign out[3468] = layer_0[4465] & ~layer_0[1392]; 
    assign out[3469] = layer_0[3347] & ~layer_0[3281]; 
    assign out[3470] = ~(layer_0[6276] & layer_0[79]); 
    assign out[3471] = ~(layer_0[5980] ^ layer_0[7718]); 
    assign out[3472] = layer_0[1247]; 
    assign out[3473] = layer_0[4073]; 
    assign out[3474] = layer_0[3300] ^ layer_0[748]; 
    assign out[3475] = ~(layer_0[2263] | layer_0[7495]); 
    assign out[3476] = layer_0[244] | layer_0[3148]; 
    assign out[3477] = ~(layer_0[6359] ^ layer_0[5336]); 
    assign out[3478] = ~(layer_0[4921] ^ layer_0[886]); 
    assign out[3479] = ~(layer_0[1642] ^ layer_0[520]); 
    assign out[3480] = ~layer_0[7226] | (layer_0[7226] & layer_0[3425]); 
    assign out[3481] = ~(layer_0[430] & layer_0[3294]); 
    assign out[3482] = layer_0[5841]; 
    assign out[3483] = ~(layer_0[7262] ^ layer_0[4961]); 
    assign out[3484] = layer_0[5515] ^ layer_0[4455]; 
    assign out[3485] = layer_0[923] ^ layer_0[5102]; 
    assign out[3486] = ~layer_0[1379] | (layer_0[1379] & layer_0[1075]); 
    assign out[3487] = layer_0[4236] ^ layer_0[5039]; 
    assign out[3488] = layer_0[270] ^ layer_0[7284]; 
    assign out[3489] = layer_0[3019] ^ layer_0[3324]; 
    assign out[3490] = ~layer_0[6075]; 
    assign out[3491] = layer_0[7219] ^ layer_0[1423]; 
    assign out[3492] = layer_0[4529]; 
    assign out[3493] = layer_0[3578] & ~layer_0[4299]; 
    assign out[3494] = layer_0[6024] & ~layer_0[7588]; 
    assign out[3495] = ~(layer_0[3053] ^ layer_0[2942]); 
    assign out[3496] = layer_0[201] ^ layer_0[5529]; 
    assign out[3497] = ~layer_0[11]; 
    assign out[3498] = layer_0[3248] ^ layer_0[5746]; 
    assign out[3499] = ~(layer_0[2431] ^ layer_0[2356]); 
    assign out[3500] = ~(layer_0[3423] ^ layer_0[6371]); 
    assign out[3501] = layer_0[7417]; 
    assign out[3502] = layer_0[2838] & layer_0[103]; 
    assign out[3503] = ~(layer_0[3876] | layer_0[4328]); 
    assign out[3504] = ~layer_0[7691] | (layer_0[7691] & layer_0[281]); 
    assign out[3505] = ~(layer_0[1524] ^ layer_0[47]); 
    assign out[3506] = ~(layer_0[4790] ^ layer_0[7720]); 
    assign out[3507] = layer_0[6824] | layer_0[5704]; 
    assign out[3508] = layer_0[3213] | layer_0[5753]; 
    assign out[3509] = layer_0[6908] ^ layer_0[4293]; 
    assign out[3510] = ~(layer_0[6619] ^ layer_0[7466]); 
    assign out[3511] = layer_0[2428] | layer_0[178]; 
    assign out[3512] = layer_0[3605] | layer_0[3307]; 
    assign out[3513] = layer_0[5929] | layer_0[5492]; 
    assign out[3514] = layer_0[994] ^ layer_0[4811]; 
    assign out[3515] = layer_0[282] & layer_0[2861]; 
    assign out[3516] = ~layer_0[2616] | (layer_0[5163] & layer_0[2616]); 
    assign out[3517] = ~layer_0[6009]; 
    assign out[3518] = ~layer_0[108] | (layer_0[108] & layer_0[2482]); 
    assign out[3519] = layer_0[824] ^ layer_0[1134]; 
    assign out[3520] = ~(layer_0[515] ^ layer_0[5314]); 
    assign out[3521] = ~(layer_0[3471] ^ layer_0[389]); 
    assign out[3522] = layer_0[1561] ^ layer_0[878]; 
    assign out[3523] = layer_0[781] & ~layer_0[6298]; 
    assign out[3524] = ~(layer_0[1692] ^ layer_0[3309]); 
    assign out[3525] = layer_0[4983] ^ layer_0[7417]; 
    assign out[3526] = layer_0[3690] & ~layer_0[3677]; 
    assign out[3527] = ~layer_0[3771] | (layer_0[3769] & layer_0[3771]); 
    assign out[3528] = ~layer_0[4429]; 
    assign out[3529] = layer_0[7225] ^ layer_0[2761]; 
    assign out[3530] = ~layer_0[1345] | (layer_0[400] & layer_0[1345]); 
    assign out[3531] = ~(layer_0[2393] ^ layer_0[7599]); 
    assign out[3532] = layer_0[7708]; 
    assign out[3533] = ~(layer_0[1275] ^ layer_0[5965]); 
    assign out[3534] = layer_0[4824] & ~layer_0[6410]; 
    assign out[3535] = layer_0[635] & ~layer_0[3583]; 
    assign out[3536] = ~(layer_0[3139] & layer_0[3040]); 
    assign out[3537] = ~(layer_0[3408] ^ layer_0[3436]); 
    assign out[3538] = ~(layer_0[4943] ^ layer_0[1168]); 
    assign out[3539] = ~(layer_0[5924] & layer_0[718]); 
    assign out[3540] = layer_0[1601]; 
    assign out[3541] = layer_0[3820]; 
    assign out[3542] = layer_0[6843] & layer_0[774]; 
    assign out[3543] = layer_0[169] & layer_0[7821]; 
    assign out[3544] = ~(layer_0[6079] ^ layer_0[1760]); 
    assign out[3545] = layer_0[4384] ^ layer_0[7800]; 
    assign out[3546] = ~(layer_0[1072] ^ layer_0[3235]); 
    assign out[3547] = layer_0[5688] & ~layer_0[5690]; 
    assign out[3548] = layer_0[6890] ^ layer_0[981]; 
    assign out[3549] = layer_0[7469] ^ layer_0[4747]; 
    assign out[3550] = ~(layer_0[913] ^ layer_0[7985]); 
    assign out[3551] = layer_0[4541]; 
    assign out[3552] = ~(layer_0[2147] & layer_0[6791]); 
    assign out[3553] = ~layer_0[7571]; 
    assign out[3554] = layer_0[3675] ^ layer_0[5328]; 
    assign out[3555] = ~(layer_0[6851] ^ layer_0[1096]); 
    assign out[3556] = ~(layer_0[5405] ^ layer_0[4116]); 
    assign out[3557] = layer_0[2545] & ~layer_0[6346]; 
    assign out[3558] = layer_0[7270] & ~layer_0[6316]; 
    assign out[3559] = layer_0[847] ^ layer_0[5508]; 
    assign out[3560] = ~(layer_0[5486] ^ layer_0[2652]); 
    assign out[3561] = layer_0[717] | layer_0[7351]; 
    assign out[3562] = layer_0[2491] ^ layer_0[7674]; 
    assign out[3563] = ~(layer_0[4050] ^ layer_0[7552]); 
    assign out[3564] = layer_0[7535] | layer_0[31]; 
    assign out[3565] = ~(layer_0[7587] & layer_0[1941]); 
    assign out[3566] = layer_0[1740] ^ layer_0[7523]; 
    assign out[3567] = ~layer_0[609] | (layer_0[7308] & layer_0[609]); 
    assign out[3568] = layer_0[2560] ^ layer_0[1590]; 
    assign out[3569] = ~(layer_0[7746] ^ layer_0[6095]); 
    assign out[3570] = layer_0[5513]; 
    assign out[3571] = layer_0[463] ^ layer_0[551]; 
    assign out[3572] = layer_0[5904] ^ layer_0[2982]; 
    assign out[3573] = ~(layer_0[7676] & layer_0[1345]); 
    assign out[3574] = ~layer_0[2886] | (layer_0[2886] & layer_0[6495]); 
    assign out[3575] = ~(layer_0[3386] ^ layer_0[3541]); 
    assign out[3576] = layer_0[2211] ^ layer_0[7078]; 
    assign out[3577] = layer_0[811] ^ layer_0[3447]; 
    assign out[3578] = layer_0[7166] ^ layer_0[4173]; 
    assign out[3579] = ~layer_0[6260]; 
    assign out[3580] = layer_0[6885] & ~layer_0[3744]; 
    assign out[3581] = layer_0[7141]; 
    assign out[3582] = ~layer_0[7860]; 
    assign out[3583] = layer_0[4926] & layer_0[4619]; 
    assign out[3584] = layer_0[286] ^ layer_0[2325]; 
    assign out[3585] = 1'b1; 
    assign out[3586] = ~layer_0[3525] | (layer_0[3767] & layer_0[3525]); 
    assign out[3587] = ~(layer_0[2737] | layer_0[4357]); 
    assign out[3588] = ~(layer_0[6100] | layer_0[4145]); 
    assign out[3589] = layer_0[2421] ^ layer_0[3298]; 
    assign out[3590] = layer_0[2571] & ~layer_0[7741]; 
    assign out[3591] = ~(layer_0[3464] & layer_0[3099]); 
    assign out[3592] = ~(layer_0[7879] | layer_0[1442]); 
    assign out[3593] = ~(layer_0[4414] ^ layer_0[2295]); 
    assign out[3594] = layer_0[6682] ^ layer_0[7946]; 
    assign out[3595] = ~(layer_0[4794] ^ layer_0[4226]); 
    assign out[3596] = ~(layer_0[2053] ^ layer_0[6426]); 
    assign out[3597] = ~(layer_0[407] ^ layer_0[373]); 
    assign out[3598] = layer_0[6401] ^ layer_0[570]; 
    assign out[3599] = layer_0[4360] ^ layer_0[4052]; 
    assign out[3600] = ~layer_0[408]; 
    assign out[3601] = layer_0[2579] & layer_0[1936]; 
    assign out[3602] = layer_0[2254] ^ layer_0[2848]; 
    assign out[3603] = ~layer_0[2115] | (layer_0[2115] & layer_0[192]); 
    assign out[3604] = ~layer_0[7894]; 
    assign out[3605] = layer_0[5372] ^ layer_0[2858]; 
    assign out[3606] = ~(layer_0[6053] ^ layer_0[1524]); 
    assign out[3607] = layer_0[3828] & ~layer_0[3161]; 
    assign out[3608] = layer_0[3545]; 
    assign out[3609] = layer_0[4337] & ~layer_0[306]; 
    assign out[3610] = layer_0[3070] ^ layer_0[2157]; 
    assign out[3611] = layer_0[1951] | layer_0[1651]; 
    assign out[3612] = ~(layer_0[5111] ^ layer_0[281]); 
    assign out[3613] = layer_0[5516] & ~layer_0[5394]; 
    assign out[3614] = ~(layer_0[1243] | layer_0[5789]); 
    assign out[3615] = layer_0[235] & layer_0[2850]; 
    assign out[3616] = layer_0[3918]; 
    assign out[3617] = layer_0[243] | layer_0[3255]; 
    assign out[3618] = layer_0[5684]; 
    assign out[3619] = layer_0[1107] & layer_0[1266]; 
    assign out[3620] = layer_0[6448] & ~layer_0[972]; 
    assign out[3621] = ~layer_0[6059] | (layer_0[6059] & layer_0[993]); 
    assign out[3622] = layer_0[3445] & ~layer_0[4629]; 
    assign out[3623] = ~(layer_0[7307] ^ layer_0[1669]); 
    assign out[3624] = ~(layer_0[3264] ^ layer_0[3210]); 
    assign out[3625] = layer_0[4488] ^ layer_0[3270]; 
    assign out[3626] = ~layer_0[2863]; 
    assign out[3627] = ~layer_0[1953]; 
    assign out[3628] = layer_0[3904]; 
    assign out[3629] = layer_0[4428] ^ layer_0[1353]; 
    assign out[3630] = 1'b0; 
    assign out[3631] = layer_0[7960] & ~layer_0[941]; 
    assign out[3632] = layer_0[5478] & layer_0[438]; 
    assign out[3633] = layer_0[6835] & layer_0[3034]; 
    assign out[3634] = ~(layer_0[2389] | layer_0[6537]); 
    assign out[3635] = layer_0[6076] | layer_0[3348]; 
    assign out[3636] = ~layer_0[6795]; 
    assign out[3637] = ~layer_0[4343]; 
    assign out[3638] = layer_0[6983] & layer_0[4850]; 
    assign out[3639] = layer_0[143] & ~layer_0[370]; 
    assign out[3640] = layer_0[5798] & ~layer_0[4823]; 
    assign out[3641] = layer_0[4693] | layer_0[7563]; 
    assign out[3642] = ~(layer_0[7630] ^ layer_0[6380]); 
    assign out[3643] = ~(layer_0[2084] ^ layer_0[2329]); 
    assign out[3644] = layer_0[3414] ^ layer_0[4648]; 
    assign out[3645] = layer_0[679] ^ layer_0[3146]; 
    assign out[3646] = layer_0[5006] | layer_0[3087]; 
    assign out[3647] = layer_0[7405] ^ layer_0[7771]; 
    assign out[3648] = layer_0[4722] & ~layer_0[596]; 
    assign out[3649] = layer_0[2982]; 
    assign out[3650] = ~(layer_0[3641] | layer_0[1993]); 
    assign out[3651] = layer_0[1086] ^ layer_0[6166]; 
    assign out[3652] = ~layer_0[855] | (layer_0[855] & layer_0[525]); 
    assign out[3653] = layer_0[1627]; 
    assign out[3654] = ~(layer_0[76] | layer_0[4731]); 
    assign out[3655] = layer_0[5223]; 
    assign out[3656] = ~layer_0[436]; 
    assign out[3657] = layer_0[6445] & ~layer_0[1714]; 
    assign out[3658] = layer_0[3451] & layer_0[3597]; 
    assign out[3659] = ~layer_0[559] | (layer_0[559] & layer_0[6296]); 
    assign out[3660] = ~(layer_0[4807] ^ layer_0[754]); 
    assign out[3661] = layer_0[1389] & ~layer_0[2123]; 
    assign out[3662] = layer_0[2999] ^ layer_0[1464]; 
    assign out[3663] = layer_0[2735] ^ layer_0[6962]; 
    assign out[3664] = layer_0[1397] ^ layer_0[7424]; 
    assign out[3665] = layer_0[6433] & ~layer_0[2801]; 
    assign out[3666] = layer_0[6882] | layer_0[2829]; 
    assign out[3667] = layer_0[4198] & ~layer_0[593]; 
    assign out[3668] = layer_0[1487] ^ layer_0[6402]; 
    assign out[3669] = ~(layer_0[1876] ^ layer_0[4749]); 
    assign out[3670] = layer_0[6464] & ~layer_0[5850]; 
    assign out[3671] = layer_0[7858]; 
    assign out[3672] = ~(layer_0[7782] | layer_0[7553]); 
    assign out[3673] = layer_0[6904] ^ layer_0[547]; 
    assign out[3674] = ~layer_0[6348] | (layer_0[7103] & layer_0[6348]); 
    assign out[3675] = ~(layer_0[4937] | layer_0[4759]); 
    assign out[3676] = layer_0[7528] & ~layer_0[958]; 
    assign out[3677] = ~layer_0[5281]; 
    assign out[3678] = ~(layer_0[1740] ^ layer_0[3907]); 
    assign out[3679] = layer_0[5460] ^ layer_0[6024]; 
    assign out[3680] = ~(layer_0[2054] ^ layer_0[404]); 
    assign out[3681] = ~layer_0[3842] | (layer_0[3842] & layer_0[7211]); 
    assign out[3682] = ~layer_0[2217]; 
    assign out[3683] = ~(layer_0[4492] ^ layer_0[783]); 
    assign out[3684] = ~layer_0[6502]; 
    assign out[3685] = ~layer_0[3193] | (layer_0[344] & layer_0[3193]); 
    assign out[3686] = layer_0[1793] | layer_0[3329]; 
    assign out[3687] = layer_0[3527] ^ layer_0[3453]; 
    assign out[3688] = layer_0[3502] | layer_0[768]; 
    assign out[3689] = layer_0[646] & ~layer_0[3549]; 
    assign out[3690] = layer_0[7322]; 
    assign out[3691] = layer_0[5274] ^ layer_0[7791]; 
    assign out[3692] = layer_0[2400] & layer_0[3595]; 
    assign out[3693] = layer_0[2812] & ~layer_0[806]; 
    assign out[3694] = ~(layer_0[1821] ^ layer_0[3543]); 
    assign out[3695] = ~layer_0[437]; 
    assign out[3696] = ~layer_0[7062] | (layer_0[7062] & layer_0[2352]); 
    assign out[3697] = layer_0[906] & ~layer_0[3841]; 
    assign out[3698] = layer_0[2607]; 
    assign out[3699] = ~(layer_0[2394] ^ layer_0[6088]); 
    assign out[3700] = layer_0[769]; 
    assign out[3701] = layer_0[3965]; 
    assign out[3702] = layer_0[291] & ~layer_0[2176]; 
    assign out[3703] = ~(layer_0[4710] ^ layer_0[6036]); 
    assign out[3704] = ~layer_0[1979]; 
    assign out[3705] = layer_0[2020] & ~layer_0[6788]; 
    assign out[3706] = layer_0[6182] ^ layer_0[5453]; 
    assign out[3707] = layer_0[65]; 
    assign out[3708] = ~layer_0[1263]; 
    assign out[3709] = layer_0[7965] & layer_0[5876]; 
    assign out[3710] = layer_0[5812]; 
    assign out[3711] = layer_0[406] ^ layer_0[3071]; 
    assign out[3712] = layer_0[688] | layer_0[7298]; 
    assign out[3713] = layer_0[6832] & ~layer_0[820]; 
    assign out[3714] = ~layer_0[2361]; 
    assign out[3715] = ~(layer_0[1550] ^ layer_0[6577]); 
    assign out[3716] = layer_0[6130] & ~layer_0[4661]; 
    assign out[3717] = layer_0[6418] & layer_0[67]; 
    assign out[3718] = layer_0[5386] & ~layer_0[7966]; 
    assign out[3719] = layer_0[7150]; 
    assign out[3720] = layer_0[5403] & ~layer_0[5437]; 
    assign out[3721] = ~layer_0[3490]; 
    assign out[3722] = layer_0[1861] & ~layer_0[6478]; 
    assign out[3723] = layer_0[3235] ^ layer_0[4570]; 
    assign out[3724] = layer_0[5915]; 
    assign out[3725] = ~(layer_0[1839] ^ layer_0[4752]); 
    assign out[3726] = layer_0[1816] & ~layer_0[1102]; 
    assign out[3727] = layer_0[6901]; 
    assign out[3728] = layer_0[3736] & ~layer_0[1237]; 
    assign out[3729] = layer_0[7100] ^ layer_0[5957]; 
    assign out[3730] = ~(layer_0[6554] ^ layer_0[7324]); 
    assign out[3731] = ~layer_0[6468]; 
    assign out[3732] = ~(layer_0[4336] ^ layer_0[847]); 
    assign out[3733] = layer_0[1269] & ~layer_0[4308]; 
    assign out[3734] = ~(layer_0[7806] ^ layer_0[5702]); 
    assign out[3735] = layer_0[3899]; 
    assign out[3736] = layer_0[1074] ^ layer_0[7916]; 
    assign out[3737] = layer_0[1517]; 
    assign out[3738] = layer_0[3774]; 
    assign out[3739] = layer_0[6985] & layer_0[7947]; 
    assign out[3740] = ~layer_0[4383] | (layer_0[2040] & layer_0[4383]); 
    assign out[3741] = ~(layer_0[7528] ^ layer_0[1802]); 
    assign out[3742] = layer_0[7148] & ~layer_0[7336]; 
    assign out[3743] = layer_0[6640] & layer_0[2160]; 
    assign out[3744] = layer_0[57]; 
    assign out[3745] = ~layer_0[6570]; 
    assign out[3746] = layer_0[3076]; 
    assign out[3747] = ~(layer_0[48] ^ layer_0[961]); 
    assign out[3748] = layer_0[3082]; 
    assign out[3749] = layer_0[3753] & ~layer_0[4356]; 
    assign out[3750] = layer_0[5091]; 
    assign out[3751] = layer_0[3829] & layer_0[5583]; 
    assign out[3752] = layer_0[3620] & ~layer_0[661]; 
    assign out[3753] = layer_0[2715] & ~layer_0[6938]; 
    assign out[3754] = layer_0[4271] & ~layer_0[2778]; 
    assign out[3755] = ~(layer_0[2182] ^ layer_0[7851]); 
    assign out[3756] = layer_0[970] ^ layer_0[3054]; 
    assign out[3757] = layer_0[2069] ^ layer_0[6305]; 
    assign out[3758] = ~(layer_0[4583] ^ layer_0[386]); 
    assign out[3759] = layer_0[203]; 
    assign out[3760] = ~layer_0[1538] | (layer_0[1538] & layer_0[3816]); 
    assign out[3761] = ~layer_0[4185] | (layer_0[4185] & layer_0[4579]); 
    assign out[3762] = ~(layer_0[5767] ^ layer_0[5320]); 
    assign out[3763] = layer_0[446] & ~layer_0[6711]; 
    assign out[3764] = ~(layer_0[1031] | layer_0[4252]); 
    assign out[3765] = layer_0[4588] & ~layer_0[5778]; 
    assign out[3766] = layer_0[2794]; 
    assign out[3767] = layer_0[5954] ^ layer_0[1375]; 
    assign out[3768] = layer_0[7285] ^ layer_0[5827]; 
    assign out[3769] = ~(layer_0[3923] & layer_0[7752]); 
    assign out[3770] = layer_0[2429] & layer_0[4452]; 
    assign out[3771] = layer_0[6634]; 
    assign out[3772] = layer_0[7178] & ~layer_0[4645]; 
    assign out[3773] = layer_0[3319]; 
    assign out[3774] = layer_0[1414] & ~layer_0[582]; 
    assign out[3775] = layer_0[4079]; 
    assign out[3776] = layer_0[1652] & ~layer_0[7609]; 
    assign out[3777] = ~(layer_0[480] ^ layer_0[7041]); 
    assign out[3778] = ~(layer_0[1190] & layer_0[654]); 
    assign out[3779] = layer_0[314] ^ layer_0[1434]; 
    assign out[3780] = ~(layer_0[1967] | layer_0[7520]); 
    assign out[3781] = ~(layer_0[7449] ^ layer_0[7162]); 
    assign out[3782] = layer_0[1506] ^ layer_0[512]; 
    assign out[3783] = ~(layer_0[7013] ^ layer_0[4296]); 
    assign out[3784] = ~(layer_0[3125] ^ layer_0[950]); 
    assign out[3785] = ~layer_0[792] | (layer_0[7472] & layer_0[792]); 
    assign out[3786] = ~layer_0[2026] | (layer_0[2026] & layer_0[3088]); 
    assign out[3787] = layer_0[2135] ^ layer_0[7903]; 
    assign out[3788] = ~layer_0[2844]; 
    assign out[3789] = ~(layer_0[6896] ^ layer_0[3610]); 
    assign out[3790] = layer_0[2148]; 
    assign out[3791] = layer_0[5669] & layer_0[1943]; 
    assign out[3792] = layer_0[4181] ^ layer_0[3942]; 
    assign out[3793] = ~layer_0[1950] | (layer_0[1950] & layer_0[7047]); 
    assign out[3794] = layer_0[3009] ^ layer_0[6034]; 
    assign out[3795] = ~(layer_0[412] | layer_0[7518]); 
    assign out[3796] = layer_0[4832] & ~layer_0[6583]; 
    assign out[3797] = layer_0[7326] & ~layer_0[4643]; 
    assign out[3798] = layer_0[787]; 
    assign out[3799] = layer_0[3574] ^ layer_0[1869]; 
    assign out[3800] = ~(layer_0[633] | layer_0[440]); 
    assign out[3801] = layer_0[7029]; 
    assign out[3802] = layer_0[6906]; 
    assign out[3803] = layer_0[7562]; 
    assign out[3804] = layer_0[7695] & layer_0[5543]; 
    assign out[3805] = layer_0[830] & ~layer_0[1172]; 
    assign out[3806] = ~(layer_0[7228] ^ layer_0[1503]); 
    assign out[3807] = ~(layer_0[6496] ^ layer_0[798]); 
    assign out[3808] = ~(layer_0[3953] ^ layer_0[584]); 
    assign out[3809] = layer_0[3194] ^ layer_0[4474]; 
    assign out[3810] = ~layer_0[4057]; 
    assign out[3811] = layer_0[648]; 
    assign out[3812] = layer_0[3262] ^ layer_0[2481]; 
    assign out[3813] = layer_0[5723] ^ layer_0[7165]; 
    assign out[3814] = ~layer_0[5125] | (layer_0[534] & layer_0[5125]); 
    assign out[3815] = ~(layer_0[5418] ^ layer_0[2272]); 
    assign out[3816] = ~(layer_0[6102] ^ layer_0[7192]); 
    assign out[3817] = ~(layer_0[2788] ^ layer_0[4840]); 
    assign out[3818] = layer_0[5351]; 
    assign out[3819] = layer_0[3559] & layer_0[1145]; 
    assign out[3820] = ~layer_0[4665]; 
    assign out[3821] = ~(layer_0[5844] ^ layer_0[6759]); 
    assign out[3822] = ~layer_0[5880] | (layer_0[5880] & layer_0[7024]); 
    assign out[3823] = ~layer_0[1809]; 
    assign out[3824] = layer_0[6362] ^ layer_0[4947]; 
    assign out[3825] = layer_0[779] & layer_0[4694]; 
    assign out[3826] = layer_0[4335] & ~layer_0[7171]; 
    assign out[3827] = layer_0[6220]; 
    assign out[3828] = ~layer_0[1011]; 
    assign out[3829] = ~(layer_0[4509] & layer_0[6080]); 
    assign out[3830] = ~layer_0[643]; 
    assign out[3831] = layer_0[6675] | layer_0[5156]; 
    assign out[3832] = layer_0[7976] ^ layer_0[4601]; 
    assign out[3833] = layer_0[14] & ~layer_0[7801]; 
    assign out[3834] = ~(layer_0[6517] ^ layer_0[3411]); 
    assign out[3835] = layer_0[6476] ^ layer_0[5546]; 
    assign out[3836] = layer_0[7131] ^ layer_0[2434]; 
    assign out[3837] = layer_0[1663]; 
    assign out[3838] = layer_0[5857] & ~layer_0[4245]; 
    assign out[3839] = ~layer_0[6335]; 
    assign out[3840] = layer_0[4235] & ~layer_0[6756]; 
    assign out[3841] = layer_0[7267] & layer_0[1473]; 
    assign out[3842] = layer_0[5489] & ~layer_0[7764]; 
    assign out[3843] = ~layer_0[1020]; 
    assign out[3844] = ~(layer_0[5363] ^ layer_0[4211]); 
    assign out[3845] = layer_0[4395] ^ layer_0[6205]; 
    assign out[3846] = layer_0[5694] ^ layer_0[3337]; 
    assign out[3847] = layer_0[1537] | layer_0[1398]; 
    assign out[3848] = layer_0[5561]; 
    assign out[3849] = layer_0[6994] | layer_0[3622]; 
    assign out[3850] = layer_0[2169] ^ layer_0[2992]; 
    assign out[3851] = layer_0[5676]; 
    assign out[3852] = layer_0[1189] & ~layer_0[3643]; 
    assign out[3853] = layer_0[7690] & layer_0[4463]; 
    assign out[3854] = layer_0[275] ^ layer_0[2298]; 
    assign out[3855] = ~(layer_0[5802] ^ layer_0[7715]); 
    assign out[3856] = layer_0[3033] & ~layer_0[3811]; 
    assign out[3857] = layer_0[637] & layer_0[2089]; 
    assign out[3858] = ~(layer_0[7632] ^ layer_0[6737]); 
    assign out[3859] = layer_0[1066] ^ layer_0[3872]; 
    assign out[3860] = ~(layer_0[7018] ^ layer_0[989]); 
    assign out[3861] = layer_0[1452] & ~layer_0[4342]; 
    assign out[3862] = layer_0[4165] & ~layer_0[381]; 
    assign out[3863] = layer_0[2262] ^ layer_0[573]; 
    assign out[3864] = ~layer_0[2556] | (layer_0[2556] & layer_0[5609]); 
    assign out[3865] = ~layer_0[7975]; 
    assign out[3866] = ~(layer_0[2646] ^ layer_0[4810]); 
    assign out[3867] = layer_0[1007] & layer_0[5685]; 
    assign out[3868] = layer_0[189] & ~layer_0[5875]; 
    assign out[3869] = layer_0[3551]; 
    assign out[3870] = ~(layer_0[3835] ^ layer_0[3032]); 
    assign out[3871] = layer_0[2928] ^ layer_0[346]; 
    assign out[3872] = ~(layer_0[7700] ^ layer_0[250]); 
    assign out[3873] = ~layer_0[3440]; 
    assign out[3874] = layer_0[1018] | layer_0[2826]; 
    assign out[3875] = layer_0[4043] | layer_0[5771]; 
    assign out[3876] = layer_0[44]; 
    assign out[3877] = layer_0[2614] ^ layer_0[3065]; 
    assign out[3878] = layer_0[1641] & layer_0[7182]; 
    assign out[3879] = layer_0[5429]; 
    assign out[3880] = ~(layer_0[64] | layer_0[5696]); 
    assign out[3881] = ~(layer_0[5491] ^ layer_0[7366]); 
    assign out[3882] = ~layer_0[5437]; 
    assign out[3883] = layer_0[5061]; 
    assign out[3884] = ~(layer_0[229] ^ layer_0[3176]); 
    assign out[3885] = layer_0[755] & layer_0[6321]; 
    assign out[3886] = layer_0[5338] ^ layer_0[2920]; 
    assign out[3887] = layer_0[2142] ^ layer_0[6110]; 
    assign out[3888] = layer_0[5567] ^ layer_0[7371]; 
    assign out[3889] = ~(layer_0[6888] ^ layer_0[2629]); 
    assign out[3890] = layer_0[1226] ^ layer_0[741]; 
    assign out[3891] = ~(layer_0[6404] ^ layer_0[1631]); 
    assign out[3892] = ~(layer_0[7389] ^ layer_0[5713]); 
    assign out[3893] = layer_0[1939] & layer_0[1720]; 
    assign out[3894] = ~(layer_0[449] ^ layer_0[2190]); 
    assign out[3895] = layer_0[3966] & layer_0[6126]; 
    assign out[3896] = ~(layer_0[2539] ^ layer_0[4547]); 
    assign out[3897] = ~(layer_0[1042] & layer_0[7742]); 
    assign out[3898] = ~(layer_0[6645] | layer_0[2004]); 
    assign out[3899] = layer_0[1419] & ~layer_0[4367]; 
    assign out[3900] = layer_0[7920]; 
    assign out[3901] = layer_0[7949] & ~layer_0[5854]; 
    assign out[3902] = layer_0[179] & ~layer_0[1301]; 
    assign out[3903] = layer_0[457] ^ layer_0[1143]; 
    assign out[3904] = layer_0[502] & ~layer_0[2778]; 
    assign out[3905] = ~layer_0[3276]; 
    assign out[3906] = ~layer_0[5989] | (layer_0[6769] & layer_0[5989]); 
    assign out[3907] = ~(layer_0[5674] ^ layer_0[881]); 
    assign out[3908] = ~(layer_0[4614] ^ layer_0[4837]); 
    assign out[3909] = ~(layer_0[7144] ^ layer_0[5389]); 
    assign out[3910] = layer_0[3116]; 
    assign out[3911] = layer_0[4035]; 
    assign out[3912] = ~(layer_0[6903] | layer_0[615]); 
    assign out[3913] = ~(layer_0[7505] & layer_0[4115]); 
    assign out[3914] = layer_0[1563] & ~layer_0[6944]; 
    assign out[3915] = ~layer_0[1508]; 
    assign out[3916] = layer_0[4831]; 
    assign out[3917] = layer_0[7754]; 
    assign out[3918] = ~(layer_0[4111] | layer_0[6749]); 
    assign out[3919] = ~(layer_0[5303] ^ layer_0[3317]); 
    assign out[3920] = layer_0[4954] ^ layer_0[410]; 
    assign out[3921] = ~(layer_0[7949] ^ layer_0[7482]); 
    assign out[3922] = layer_0[1606] & ~layer_0[7438]; 
    assign out[3923] = layer_0[4975] & layer_0[2931]; 
    assign out[3924] = ~layer_0[5762]; 
    assign out[3925] = layer_0[2391] ^ layer_0[1589]; 
    assign out[3926] = ~(layer_0[1713] ^ layer_0[3647]); 
    assign out[3927] = layer_0[3008] ^ layer_0[3566]; 
    assign out[3928] = layer_0[2651]; 
    assign out[3929] = ~layer_0[1260]; 
    assign out[3930] = ~layer_0[5944]; 
    assign out[3931] = ~layer_0[2908]; 
    assign out[3932] = ~layer_0[2205]; 
    assign out[3933] = layer_0[200]; 
    assign out[3934] = layer_0[1552] & layer_0[6267]; 
    assign out[3935] = ~(layer_0[5518] ^ layer_0[5883]); 
    assign out[3936] = layer_0[3449] & ~layer_0[5571]; 
    assign out[3937] = layer_0[3804] ^ layer_0[5483]; 
    assign out[3938] = layer_0[7881] & ~layer_0[2013]; 
    assign out[3939] = layer_0[2695]; 
    assign out[3940] = layer_0[5725]; 
    assign out[3941] = ~(layer_0[2548] ^ layer_0[3211]); 
    assign out[3942] = layer_0[6221] ^ layer_0[7227]; 
    assign out[3943] = layer_0[2594] ^ layer_0[3816]; 
    assign out[3944] = ~layer_0[1299]; 
    assign out[3945] = ~(layer_0[1557] ^ layer_0[6692]); 
    assign out[3946] = layer_0[6480] & ~layer_0[1026]; 
    assign out[3947] = ~layer_0[3798]; 
    assign out[3948] = ~layer_0[7497] | (layer_0[7497] & layer_0[6143]); 
    assign out[3949] = ~layer_0[5213]; 
    assign out[3950] = layer_0[5681]; 
    assign out[3951] = ~(layer_0[577] ^ layer_0[5189]); 
    assign out[3952] = ~layer_0[1236]; 
    assign out[3953] = ~(layer_0[2688] & layer_0[475]); 
    assign out[3954] = layer_0[2109] & layer_0[4758]; 
    assign out[3955] = ~(layer_0[4553] ^ layer_0[4622]); 
    assign out[3956] = layer_0[5309] & ~layer_0[7493]; 
    assign out[3957] = layer_0[4591] & ~layer_0[7026]; 
    assign out[3958] = layer_0[2881] & layer_0[3220]; 
    assign out[3959] = ~(layer_0[6342] ^ layer_0[5252]); 
    assign out[3960] = layer_0[3776] ^ layer_0[4029]; 
    assign out[3961] = ~layer_0[545]; 
    assign out[3962] = ~layer_0[6243]; 
    assign out[3963] = layer_0[6155]; 
    assign out[3964] = layer_0[5325] & layer_0[7423]; 
    assign out[3965] = layer_0[5865]; 
    assign out[3966] = ~(layer_0[4450] | layer_0[5895]); 
    assign out[3967] = layer_0[2186] & layer_0[4325]; 
    assign out[3968] = layer_0[2056] & layer_0[3483]; 
    assign out[3969] = ~layer_0[4514] | (layer_0[4514] & layer_0[1914]); 
    assign out[3970] = ~layer_0[6235] | (layer_0[6235] & layer_0[6710]); 
    assign out[3971] = layer_0[5974] | layer_0[3733]; 
    assign out[3972] = layer_0[5172] & ~layer_0[3743]; 
    assign out[3973] = layer_0[2742]; 
    assign out[3974] = layer_0[3313] & ~layer_0[6555]; 
    assign out[3975] = ~(layer_0[5102] ^ layer_0[5151]); 
    assign out[3976] = ~layer_0[2238]; 
    assign out[3977] = layer_0[4793] & layer_0[2315]; 
    assign out[3978] = layer_0[4389] & layer_0[3656]; 
    assign out[3979] = layer_0[5085] ^ layer_0[2045]; 
    assign out[3980] = layer_0[1060] ^ layer_0[1973]; 
    assign out[3981] = layer_0[1300] & layer_0[4873]; 
    assign out[3982] = ~(layer_0[4088] & layer_0[1280]); 
    assign out[3983] = layer_0[3784] ^ layer_0[2033]; 
    assign out[3984] = ~layer_0[503]; 
    assign out[3985] = layer_0[4303] & ~layer_0[7382]; 
    assign out[3986] = layer_0[1499] ^ layer_0[2658]; 
    assign out[3987] = ~layer_0[24]; 
    assign out[3988] = ~layer_0[3081] | (layer_0[2892] & layer_0[3081]); 
    assign out[3989] = ~(layer_0[931] | layer_0[5574]); 
    assign out[3990] = layer_0[7186]; 
    assign out[3991] = layer_0[3649] & ~layer_0[7228]; 
    assign out[3992] = layer_0[7160] & ~layer_0[4218]; 
    assign out[3993] = layer_0[7855] & ~layer_0[7196]; 
    assign out[3994] = layer_0[7862] ^ layer_0[4655]; 
    assign out[3995] = ~layer_0[7596]; 
    assign out[3996] = ~(layer_0[2754] ^ layer_0[4662]); 
    assign out[3997] = layer_0[5328] & ~layer_0[5520]; 
    assign out[3998] = ~layer_0[1103] | (layer_0[5041] & layer_0[1103]); 
    assign out[3999] = ~(layer_0[401] ^ layer_0[5187]); 
    assign out[4000] = layer_0[7328] ^ layer_0[294]; 
    assign out[4001] = layer_0[4922]; 
    assign out[4002] = layer_0[4262] ^ layer_0[2083]; 
    assign out[4003] = ~layer_0[1271] | (layer_0[1271] & layer_0[5232]); 
    assign out[4004] = layer_0[7729] ^ layer_0[7142]; 
    assign out[4005] = ~layer_0[669]; 
    assign out[4006] = layer_0[2152]; 
    assign out[4007] = ~(layer_0[7554] & layer_0[1576]); 
    assign out[4008] = ~(layer_0[4647] & layer_0[6819]); 
    assign out[4009] = ~(layer_0[3921] ^ layer_0[4722]); 
    assign out[4010] = layer_0[5839]; 
    assign out[4011] = ~(layer_0[6113] | layer_0[2233]); 
    assign out[4012] = ~(layer_0[836] & layer_0[3783]); 
    assign out[4013] = layer_0[6082] & ~layer_0[6530]; 
    assign out[4014] = ~layer_0[3410]; 
    assign out[4015] = ~(layer_0[1832] ^ layer_0[5627]); 
    assign out[4016] = ~layer_0[6297] | (layer_0[6297] & layer_0[553]); 
    assign out[4017] = layer_0[1448]; 
    assign out[4018] = layer_0[3630]; 
    assign out[4019] = layer_0[6455] & ~layer_0[360]; 
    assign out[4020] = ~layer_0[3666] | (layer_0[4241] & layer_0[3666]); 
    assign out[4021] = layer_0[6811] ^ layer_0[1708]; 
    assign out[4022] = layer_0[3621]; 
    assign out[4023] = layer_0[799] & ~layer_0[4890]; 
    assign out[4024] = layer_0[7731] & ~layer_0[3571]; 
    assign out[4025] = ~layer_0[357] | (layer_0[2268] & layer_0[357]); 
    assign out[4026] = layer_0[7043]; 
    assign out[4027] = layer_0[6652] ^ layer_0[5796]; 
    assign out[4028] = ~(layer_0[3260] ^ layer_0[640]); 
    assign out[4029] = ~(layer_0[6304] ^ layer_0[2601]); 
    assign out[4030] = layer_0[6280] ^ layer_0[3221]; 
    assign out[4031] = layer_0[5567] & ~layer_0[7756]; 
    assign out[4032] = ~(layer_0[4398] ^ layer_0[1541]); 
    assign out[4033] = layer_0[7837] ^ layer_0[739]; 
    assign out[4034] = layer_0[2255] ^ layer_0[6927]; 
    assign out[4035] = ~(layer_0[5387] & layer_0[2204]); 
    assign out[4036] = ~(layer_0[7107] ^ layer_0[3960]); 
    assign out[4037] = layer_0[3075] & ~layer_0[3428]; 
    assign out[4038] = layer_0[2981] ^ layer_0[7959]; 
    assign out[4039] = layer_0[6256] & layer_0[5449]; 
    assign out[4040] = ~layer_0[7471]; 
    assign out[4041] = ~layer_0[4512]; 
    assign out[4042] = layer_0[242] | layer_0[7287]; 
    assign out[4043] = ~(layer_0[182] ^ layer_0[7436]); 
    assign out[4044] = layer_0[1049]; 
    assign out[4045] = 1'b0; 
    assign out[4046] = ~layer_0[4427]; 
    assign out[4047] = layer_0[6501]; 
    assign out[4048] = layer_0[2481] & ~layer_0[4892]; 
    assign out[4049] = ~(layer_0[5153] & layer_0[2246]); 
    assign out[4050] = ~(layer_0[3530] ^ layer_0[2223]); 
    assign out[4051] = layer_0[1622]; 
    assign out[4052] = layer_0[4874] & ~layer_0[2435]; 
    assign out[4053] = ~(layer_0[3671] ^ layer_0[4290]); 
    assign out[4054] = layer_0[4603]; 
    assign out[4055] = layer_0[4716] ^ layer_0[6443]; 
    assign out[4056] = ~(layer_0[2224] ^ layer_0[1]); 
    assign out[4057] = layer_0[2282] & layer_0[7611]; 
    assign out[4058] = layer_0[7614]; 
    assign out[4059] = layer_0[2209]; 
    assign out[4060] = ~layer_0[1412]; 
    assign out[4061] = layer_0[4032] ^ layer_0[2903]; 
    assign out[4062] = ~(layer_0[6757] | layer_0[5711]); 
    assign out[4063] = layer_0[2422]; 
    assign out[4064] = ~(layer_0[4232] | layer_0[3258]); 
    assign out[4065] = layer_0[6531] | layer_0[7332]; 
    assign out[4066] = ~(layer_0[1971] ^ layer_0[1294]); 
    assign out[4067] = ~(layer_0[3168] ^ layer_0[1830]); 
    assign out[4068] = layer_0[4498]; 
    assign out[4069] = layer_0[1418] & ~layer_0[1099]; 
    assign out[4070] = layer_0[3910] & layer_0[2419]; 
    assign out[4071] = layer_0[871] & ~layer_0[596]; 
    assign out[4072] = ~layer_0[7634]; 
    assign out[4073] = ~layer_0[2344]; 
    assign out[4074] = ~layer_0[479]; 
    assign out[4075] = ~(layer_0[1335] | layer_0[4419]); 
    assign out[4076] = ~layer_0[1555]; 
    assign out[4077] = layer_0[6721] & layer_0[4848]; 
    assign out[4078] = layer_0[1403] ^ layer_0[6173]; 
    assign out[4079] = layer_0[2752] ^ layer_0[217]; 
    assign out[4080] = ~(layer_0[7788] | layer_0[4160]); 
    assign out[4081] = layer_0[484] ^ layer_0[6406]; 
    assign out[4082] = layer_0[1699] & layer_0[6011]; 
    assign out[4083] = ~(layer_0[5833] ^ layer_0[6338]); 
    assign out[4084] = layer_0[7249] ^ layer_0[788]; 
    assign out[4085] = layer_0[234]; 
    assign out[4086] = layer_0[1939] & layer_0[5400]; 
    assign out[4087] = ~(layer_0[3653] | layer_0[4331]); 
    assign out[4088] = ~(layer_0[5311] ^ layer_0[2215]); 
    assign out[4089] = layer_0[3647] & ~layer_0[1603]; 
    assign out[4090] = ~layer_0[505] | (layer_0[7798] & layer_0[505]); 
    assign out[4091] = ~(layer_0[4575] ^ layer_0[6693]); 
    assign out[4092] = layer_0[2633] & layer_0[6650]; 
    assign out[4093] = layer_0[7565] ^ layer_0[7321]; 
    assign out[4094] = ~layer_0[4193]; 
    assign out[4095] = ~(layer_0[6780] ^ layer_0[964]); 
    assign out[4096] = ~(layer_0[1199] ^ layer_0[7347]); 
    assign out[4097] = layer_0[7277] ^ layer_0[3286]; 
    assign out[4098] = ~(layer_0[2057] | layer_0[4934]); 
    assign out[4099] = ~layer_0[4796] | (layer_0[4796] & layer_0[609]); 
    assign out[4100] = layer_0[4351] ^ layer_0[7368]; 
    assign out[4101] = layer_0[6479] ^ layer_0[6043]; 
    assign out[4102] = ~(layer_0[3261] ^ layer_0[7090]); 
    assign out[4103] = layer_0[5183] ^ layer_0[7221]; 
    assign out[4104] = layer_0[3784] ^ layer_0[5499]; 
    assign out[4105] = ~layer_0[1446] | (layer_0[5620] & layer_0[1446]); 
    assign out[4106] = layer_0[5442]; 
    assign out[4107] = ~(layer_0[6188] ^ layer_0[4767]); 
    assign out[4108] = ~layer_0[6657] | (layer_0[4305] & layer_0[6657]); 
    assign out[4109] = ~(layer_0[5157] ^ layer_0[1297]); 
    assign out[4110] = ~(layer_0[1194] | layer_0[4585]); 
    assign out[4111] = ~(layer_0[7775] & layer_0[5253]); 
    assign out[4112] = ~(layer_0[5147] & layer_0[3403]); 
    assign out[4113] = ~(layer_0[4612] ^ layer_0[4605]); 
    assign out[4114] = layer_0[2517] ^ layer_0[2065]; 
    assign out[4115] = layer_0[5765] & layer_0[148]; 
    assign out[4116] = ~(layer_0[5099] ^ layer_0[6764]); 
    assign out[4117] = ~(layer_0[4436] ^ layer_0[433]); 
    assign out[4118] = layer_0[1754] ^ layer_0[7235]; 
    assign out[4119] = ~(layer_0[6098] ^ layer_0[7129]); 
    assign out[4120] = layer_0[6935] ^ layer_0[2030]; 
    assign out[4121] = layer_0[7352] | layer_0[4248]; 
    assign out[4122] = layer_0[2195] ^ layer_0[249]; 
    assign out[4123] = ~(layer_0[1327] ^ layer_0[548]); 
    assign out[4124] = ~(layer_0[510] & layer_0[1638]); 
    assign out[4125] = ~(layer_0[5907] | layer_0[4137]); 
    assign out[4126] = ~layer_0[1570] | (layer_0[6702] & layer_0[1570]); 
    assign out[4127] = ~(layer_0[3204] ^ layer_0[6910]); 
    assign out[4128] = layer_0[2733]; 
    assign out[4129] = ~(layer_0[2472] ^ layer_0[7818]); 
    assign out[4130] = layer_0[5469] | layer_0[2462]; 
    assign out[4131] = layer_0[6240] & layer_0[6269]; 
    assign out[4132] = ~(layer_0[5330] ^ layer_0[7392]); 
    assign out[4133] = layer_0[2101] ^ layer_0[3859]; 
    assign out[4134] = layer_0[7102] ^ layer_0[1037]; 
    assign out[4135] = ~(layer_0[5795] ^ layer_0[1008]); 
    assign out[4136] = ~layer_0[7130] | (layer_0[7130] & layer_0[1839]); 
    assign out[4137] = layer_0[6565] ^ layer_0[2186]; 
    assign out[4138] = layer_0[4437] ^ layer_0[3154]; 
    assign out[4139] = layer_0[7156] ^ layer_0[2732]; 
    assign out[4140] = ~(layer_0[5419] ^ layer_0[4081]); 
    assign out[4141] = layer_0[7880]; 
    assign out[4142] = layer_0[185] ^ layer_0[1731]; 
    assign out[4143] = layer_0[6223] ^ layer_0[223]; 
    assign out[4144] = ~layer_0[3538] | (layer_0[7479] & layer_0[3538]); 
    assign out[4145] = layer_0[6219] & ~layer_0[603]; 
    assign out[4146] = layer_0[1361] | layer_0[5056]; 
    assign out[4147] = ~layer_0[7313]; 
    assign out[4148] = ~(layer_0[3780] & layer_0[1447]); 
    assign out[4149] = layer_0[6055] ^ layer_0[6719]; 
    assign out[4150] = ~layer_0[2522]; 
    assign out[4151] = ~(layer_0[7645] ^ layer_0[6602]); 
    assign out[4152] = layer_0[6163] & ~layer_0[5576]; 
    assign out[4153] = layer_0[4588] ^ layer_0[3694]; 
    assign out[4154] = ~layer_0[6408] | (layer_0[1382] & layer_0[6408]); 
    assign out[4155] = layer_0[5192] ^ layer_0[6233]; 
    assign out[4156] = layer_0[5272] ^ layer_0[3994]; 
    assign out[4157] = ~(layer_0[7654] ^ layer_0[295]); 
    assign out[4158] = ~layer_0[132]; 
    assign out[4159] = ~layer_0[7128] | (layer_0[7128] & layer_0[5856]); 
    assign out[4160] = ~(layer_0[3268] ^ layer_0[7591]); 
    assign out[4161] = ~(layer_0[383] & layer_0[574]); 
    assign out[4162] = ~(layer_0[1295] ^ layer_0[7054]); 
    assign out[4163] = layer_0[7371] ^ layer_0[6976]; 
    assign out[4164] = ~(layer_0[267] & layer_0[4077]); 
    assign out[4165] = ~(layer_0[1856] ^ layer_0[7038]); 
    assign out[4166] = ~(layer_0[7197] ^ layer_0[771]); 
    assign out[4167] = layer_0[7299] ^ layer_0[1096]; 
    assign out[4168] = ~layer_0[7714] | (layer_0[7714] & layer_0[3850]); 
    assign out[4169] = layer_0[6099] & ~layer_0[7757]; 
    assign out[4170] = layer_0[2698] ^ layer_0[4770]; 
    assign out[4171] = ~layer_0[2927] | (layer_0[4503] & layer_0[2927]); 
    assign out[4172] = ~layer_0[6922]; 
    assign out[4173] = layer_0[3952] ^ layer_0[726]; 
    assign out[4174] = layer_0[2334] | layer_0[711]; 
    assign out[4175] = ~(layer_0[5294] & layer_0[360]); 
    assign out[4176] = ~layer_0[3818]; 
    assign out[4177] = layer_0[1082] & layer_0[6007]; 
    assign out[4178] = ~layer_0[109] | (layer_0[109] & layer_0[2766]); 
    assign out[4179] = ~layer_0[7504]; 
    assign out[4180] = ~(layer_0[6177] ^ layer_0[3845]); 
    assign out[4181] = layer_0[4777] ^ layer_0[4908]; 
    assign out[4182] = layer_0[3230] & ~layer_0[5612]; 
    assign out[4183] = ~layer_0[6967] | (layer_0[3318] & layer_0[6967]); 
    assign out[4184] = ~layer_0[6285]; 
    assign out[4185] = layer_0[2337]; 
    assign out[4186] = ~(layer_0[3812] ^ layer_0[813]); 
    assign out[4187] = layer_0[2599] ^ layer_0[7059]; 
    assign out[4188] = ~(layer_0[7922] ^ layer_0[1813]); 
    assign out[4189] = layer_0[1964] & ~layer_0[6919]; 
    assign out[4190] = ~layer_0[3875] | (layer_0[3875] & layer_0[7067]); 
    assign out[4191] = layer_0[7413]; 
    assign out[4192] = layer_0[4056] | layer_0[541]; 
    assign out[4193] = layer_0[1764] ^ layer_0[1367]; 
    assign out[4194] = ~(layer_0[7857] | layer_0[6336]); 
    assign out[4195] = ~layer_0[7577]; 
    assign out[4196] = ~(layer_0[1850] | layer_0[5933]); 
    assign out[4197] = ~layer_0[7939]; 
    assign out[4198] = layer_0[6216] ^ layer_0[164]; 
    assign out[4199] = layer_0[5541] ^ layer_0[3393]; 
    assign out[4200] = layer_0[5306]; 
    assign out[4201] = layer_0[1855] | layer_0[2590]; 
    assign out[4202] = ~(layer_0[2851] ^ layer_0[2830]); 
    assign out[4203] = ~(layer_0[4834] & layer_0[1750]); 
    assign out[4204] = layer_0[5201]; 
    assign out[4205] = ~(layer_0[597] ^ layer_0[4413]); 
    assign out[4206] = layer_0[3834]; 
    assign out[4207] = layer_0[2639]; 
    assign out[4208] = ~(layer_0[2543] ^ layer_0[2543]); 
    assign out[4209] = ~layer_0[2399]; 
    assign out[4210] = ~layer_0[300]; 
    assign out[4211] = layer_0[4093]; 
    assign out[4212] = layer_0[1737] ^ layer_0[1505]; 
    assign out[4213] = ~layer_0[1128] | (layer_0[1128] & layer_0[2759]); 
    assign out[4214] = ~(layer_0[7268] ^ layer_0[3206]); 
    assign out[4215] = ~(layer_0[1787] ^ layer_0[1470]); 
    assign out[4216] = layer_0[2600] ^ layer_0[694]; 
    assign out[4217] = ~layer_0[3940] | (layer_0[3940] & layer_0[6347]); 
    assign out[4218] = ~layer_0[1984] | (layer_0[1360] & layer_0[1984]); 
    assign out[4219] = layer_0[6345] & layer_0[7066]; 
    assign out[4220] = layer_0[2231] | layer_0[3228]; 
    assign out[4221] = layer_0[1222] ^ layer_0[5017]; 
    assign out[4222] = ~layer_0[3039]; 
    assign out[4223] = ~(layer_0[3084] & layer_0[2821]); 
    assign out[4224] = layer_0[5196] ^ layer_0[2897]; 
    assign out[4225] = ~layer_0[3488] | (layer_0[3488] & layer_0[5055]); 
    assign out[4226] = ~(layer_0[4406] ^ layer_0[905]); 
    assign out[4227] = ~(layer_0[2608] ^ layer_0[5760]); 
    assign out[4228] = ~(layer_0[552] ^ layer_0[4678]); 
    assign out[4229] = ~(layer_0[5884] & layer_0[2252]); 
    assign out[4230] = ~layer_0[823]; 
    assign out[4231] = layer_0[7958] ^ layer_0[5155]; 
    assign out[4232] = layer_0[4094] & ~layer_0[990]; 
    assign out[4233] = layer_0[145] ^ layer_0[6931]; 
    assign out[4234] = layer_0[6475] ^ layer_0[5572]; 
    assign out[4235] = layer_0[3586] | layer_0[1083]; 
    assign out[4236] = layer_0[2798] ^ layer_0[5163]; 
    assign out[4237] = ~layer_0[7354] | (layer_0[5887] & layer_0[7354]); 
    assign out[4238] = layer_0[4451] ^ layer_0[3302]; 
    assign out[4239] = layer_0[2009] & layer_0[794]; 
    assign out[4240] = layer_0[2077] ^ layer_0[6807]; 
    assign out[4241] = ~(layer_0[2720] ^ layer_0[4732]); 
    assign out[4242] = layer_0[93] ^ layer_0[4289]; 
    assign out[4243] = ~(layer_0[7517] & layer_0[3300]); 
    assign out[4244] = ~(layer_0[2541] ^ layer_0[681]); 
    assign out[4245] = layer_0[3172]; 
    assign out[4246] = ~(layer_0[1600] & layer_0[1209]); 
    assign out[4247] = layer_0[7869]; 
    assign out[4248] = layer_0[2976] ^ layer_0[5175]; 
    assign out[4249] = layer_0[3328] ^ layer_0[7693]; 
    assign out[4250] = ~layer_0[1808]; 
    assign out[4251] = ~(layer_0[3237] ^ layer_0[7272]); 
    assign out[4252] = ~layer_0[1957] | (layer_0[2913] & layer_0[1957]); 
    assign out[4253] = ~layer_0[948] | (layer_0[948] & layer_0[738]); 
    assign out[4254] = layer_0[7882]; 
    assign out[4255] = layer_0[4364]; 
    assign out[4256] = ~(layer_0[7314] ^ layer_0[4328]); 
    assign out[4257] = ~(layer_0[5851] ^ layer_0[1501]); 
    assign out[4258] = ~layer_0[4240]; 
    assign out[4259] = layer_0[2284] | layer_0[1123]; 
    assign out[4260] = layer_0[6632] ^ layer_0[7928]; 
    assign out[4261] = layer_0[2642] | layer_0[2203]; 
    assign out[4262] = layer_0[750]; 
    assign out[4263] = layer_0[4070] ^ layer_0[797]; 
    assign out[4264] = ~(layer_0[7265] ^ layer_0[5230]); 
    assign out[4265] = ~(layer_0[1278] ^ layer_0[2494]); 
    assign out[4266] = ~layer_0[1566]; 
    assign out[4267] = layer_0[4269]; 
    assign out[4268] = ~(layer_0[5315] | layer_0[3866]); 
    assign out[4269] = ~layer_0[4668] | (layer_0[1439] & layer_0[4668]); 
    assign out[4270] = layer_0[3814]; 
    assign out[4271] = ~(layer_0[4768] ^ layer_0[2687]); 
    assign out[4272] = ~(layer_0[1769] ^ layer_0[4951]); 
    assign out[4273] = layer_0[3375] | layer_0[2355]; 
    assign out[4274] = ~layer_0[4367] | (layer_0[4367] & layer_0[5650]); 
    assign out[4275] = ~(layer_0[7637] ^ layer_0[7780]); 
    assign out[4276] = ~layer_0[683]; 
    assign out[4277] = ~(layer_0[5748] ^ layer_0[3862]); 
    assign out[4278] = ~layer_0[3642] | (layer_0[3642] & layer_0[3980]); 
    assign out[4279] = ~(layer_0[6337] ^ layer_0[5547]); 
    assign out[4280] = layer_0[1900] & ~layer_0[1840]; 
    assign out[4281] = layer_0[6895] | layer_0[2990]; 
    assign out[4282] = ~layer_0[2407] | (layer_0[2407] & layer_0[2068]); 
    assign out[4283] = ~layer_0[6040]; 
    assign out[4284] = ~layer_0[491] | (layer_0[6611] & layer_0[491]); 
    assign out[4285] = layer_0[167] ^ layer_0[5706]; 
    assign out[4286] = layer_0[7210] ^ layer_0[2172]; 
    assign out[4287] = layer_0[2694] ^ layer_0[6608]; 
    assign out[4288] = ~layer_0[2937] | (layer_0[1257] & layer_0[2937]); 
    assign out[4289] = layer_0[7651] | layer_0[3646]; 
    assign out[4290] = ~layer_0[868] | (layer_0[7816] & layer_0[868]); 
    assign out[4291] = layer_0[2832]; 
    assign out[4292] = layer_0[5919] ^ layer_0[839]; 
    assign out[4293] = ~(layer_0[7163] ^ layer_0[6390]); 
    assign out[4294] = layer_0[3757]; 
    assign out[4295] = ~(layer_0[2312] | layer_0[2895]); 
    assign out[4296] = layer_0[4972]; 
    assign out[4297] = ~(layer_0[2455] ^ layer_0[6078]); 
    assign out[4298] = ~layer_0[1969] | (layer_0[4536] & layer_0[1969]); 
    assign out[4299] = ~layer_0[1777]; 
    assign out[4300] = ~layer_0[5015]; 
    assign out[4301] = ~(layer_0[6172] ^ layer_0[2365]); 
    assign out[4302] = ~layer_0[1768] | (layer_0[1768] & layer_0[7572]); 
    assign out[4303] = layer_0[1205] ^ layer_0[2705]; 
    assign out[4304] = layer_0[6642] ^ layer_0[120]; 
    assign out[4305] = ~(layer_0[3316] ^ layer_0[2390]); 
    assign out[4306] = ~(layer_0[1612] ^ layer_0[3863]); 
    assign out[4307] = ~layer_0[4714]; 
    assign out[4308] = ~layer_0[1285] | (layer_0[1285] & layer_0[3350]); 
    assign out[4309] = ~(layer_0[2395] ^ layer_0[3537]); 
    assign out[4310] = layer_0[5184]; 
    assign out[4311] = ~layer_0[7890] | (layer_0[5860] & layer_0[7890]); 
    assign out[4312] = layer_0[1614] ^ layer_0[2729]; 
    assign out[4313] = ~layer_0[4647]; 
    assign out[4314] = ~layer_0[2024] | (layer_0[2024] & layer_0[3059]); 
    assign out[4315] = ~layer_0[2680]; 
    assign out[4316] = ~layer_0[5590] | (layer_0[4839] & layer_0[5590]); 
    assign out[4317] = layer_0[1230] ^ layer_0[563]; 
    assign out[4318] = ~(layer_0[7496] ^ layer_0[6042]); 
    assign out[4319] = layer_0[6401] ^ layer_0[72]; 
    assign out[4320] = layer_0[841] ^ layer_0[6894]; 
    assign out[4321] = ~layer_0[6403]; 
    assign out[4322] = ~layer_0[4151]; 
    assign out[4323] = layer_0[7953]; 
    assign out[4324] = layer_0[6336] ^ layer_0[3854]; 
    assign out[4325] = ~layer_0[6723]; 
    assign out[4326] = ~layer_0[43]; 
    assign out[4327] = layer_0[1842] ^ layer_0[2120]; 
    assign out[4328] = ~(layer_0[780] ^ layer_0[7240]); 
    assign out[4329] = layer_0[1006]; 
    assign out[4330] = ~(layer_0[3251] & layer_0[2871]); 
    assign out[4331] = layer_0[3367] ^ layer_0[1129]; 
    assign out[4332] = ~layer_0[5454]; 
    assign out[4333] = ~(layer_0[5064] ^ layer_0[979]); 
    assign out[4334] = layer_0[334]; 
    assign out[4335] = ~(layer_0[1084] ^ layer_0[1906]); 
    assign out[4336] = layer_0[5650]; 
    assign out[4337] = ~layer_0[2274] | (layer_0[2274] & layer_0[6476]); 
    assign out[4338] = layer_0[5304] | layer_0[3376]; 
    assign out[4339] = layer_0[1797] ^ layer_0[7973]; 
    assign out[4340] = layer_0[3102] ^ layer_0[6013]; 
    assign out[4341] = ~(layer_0[1691] & layer_0[2085]); 
    assign out[4342] = layer_0[4387] ^ layer_0[268]; 
    assign out[4343] = ~(layer_0[4527] ^ layer_0[1779]); 
    assign out[4344] = ~layer_0[2576]; 
    assign out[4345] = ~layer_0[1861] | (layer_0[1861] & layer_0[5194]); 
    assign out[4346] = ~layer_0[7392] | (layer_0[7792] & layer_0[7392]); 
    assign out[4347] = layer_0[2317] ^ layer_0[5358]; 
    assign out[4348] = layer_0[5819] & layer_0[1250]; 
    assign out[4349] = ~(layer_0[6272] | layer_0[5821]); 
    assign out[4350] = layer_0[394] & ~layer_0[7231]; 
    assign out[4351] = layer_0[6324] & ~layer_0[689]; 
    assign out[4352] = layer_0[2139] & ~layer_0[5530]; 
    assign out[4353] = layer_0[4521] ^ layer_0[6738]; 
    assign out[4354] = ~(layer_0[4867] & layer_0[2110]); 
    assign out[4355] = layer_0[6018] ^ layer_0[3612]; 
    assign out[4356] = ~layer_0[4092]; 
    assign out[4357] = layer_0[6131]; 
    assign out[4358] = ~(layer_0[3393] | layer_0[5196]); 
    assign out[4359] = layer_0[7411]; 
    assign out[4360] = ~(layer_0[1161] & layer_0[6397]); 
    assign out[4361] = layer_0[7167] & layer_0[4266]; 
    assign out[4362] = ~(layer_0[7152] ^ layer_0[7765]); 
    assign out[4363] = layer_0[2247]; 
    assign out[4364] = ~(layer_0[7484] ^ layer_0[5768]); 
    assign out[4365] = layer_0[7399] ^ layer_0[4998]; 
    assign out[4366] = layer_0[5264] | layer_0[3930]; 
    assign out[4367] = ~(layer_0[6926] ^ layer_0[327]); 
    assign out[4368] = layer_0[6742] ^ layer_0[3981]; 
    assign out[4369] = layer_0[1169] ^ layer_0[1548]; 
    assign out[4370] = layer_0[6525] & layer_0[2082]; 
    assign out[4371] = layer_0[3598] ^ layer_0[879]; 
    assign out[4372] = layer_0[1551]; 
    assign out[4373] = ~layer_0[5937] | (layer_0[1959] & layer_0[5937]); 
    assign out[4374] = layer_0[3978] & ~layer_0[814]; 
    assign out[4375] = ~(layer_0[3596] ^ layer_0[3883]); 
    assign out[4376] = ~(layer_0[1795] ^ layer_0[5288]); 
    assign out[4377] = ~(layer_0[7368] ^ layer_0[5235]); 
    assign out[4378] = ~(layer_0[2813] & layer_0[3844]); 
    assign out[4379] = layer_0[7018] ^ layer_0[6961]; 
    assign out[4380] = layer_0[7766] | layer_0[3619]; 
    assign out[4381] = ~layer_0[2572] | (layer_0[6884] & layer_0[2572]); 
    assign out[4382] = ~(layer_0[7452] ^ layer_0[7064]); 
    assign out[4383] = ~layer_0[453]; 
    assign out[4384] = ~layer_0[7271]; 
    assign out[4385] = layer_0[3]; 
    assign out[4386] = ~(layer_0[4434] & layer_0[4495]); 
    assign out[4387] = ~layer_0[5589]; 
    assign out[4388] = layer_0[1709] ^ layer_0[3727]; 
    assign out[4389] = ~(layer_0[5712] & layer_0[7801]); 
    assign out[4390] = layer_0[55]; 
    assign out[4391] = layer_0[6455] ^ layer_0[4462]; 
    assign out[4392] = layer_0[7349] ^ layer_0[4673]; 
    assign out[4393] = ~(layer_0[1655] | layer_0[2383]); 
    assign out[4394] = ~(layer_0[2441] ^ layer_0[3141]); 
    assign out[4395] = layer_0[5081] ^ layer_0[3649]; 
    assign out[4396] = ~(layer_0[265] & layer_0[2539]); 
    assign out[4397] = layer_0[3305] ^ layer_0[317]; 
    assign out[4398] = ~layer_0[4568]; 
    assign out[4399] = ~layer_0[5028]; 
    assign out[4400] = ~layer_0[506] | (layer_0[1101] & layer_0[506]); 
    assign out[4401] = ~layer_0[4797]; 
    assign out[4402] = layer_0[3577]; 
    assign out[4403] = ~(layer_0[7310] & layer_0[3444]); 
    assign out[4404] = layer_0[2520] & layer_0[5616]; 
    assign out[4405] = ~(layer_0[6017] & layer_0[758]); 
    assign out[4406] = layer_0[6194] ^ layer_0[6981]; 
    assign out[4407] = ~layer_0[5999]; 
    assign out[4408] = layer_0[6493] ^ layer_0[3638]; 
    assign out[4409] = layer_0[741] ^ layer_0[99]; 
    assign out[4410] = ~layer_0[5805]; 
    assign out[4411] = layer_0[5064] & layer_0[665]; 
    assign out[4412] = ~layer_0[1890]; 
    assign out[4413] = layer_0[5332] ^ layer_0[3701]; 
    assign out[4414] = layer_0[2452]; 
    assign out[4415] = ~layer_0[5261] | (layer_0[6929] & layer_0[5261]); 
    assign out[4416] = layer_0[3261] ^ layer_0[2106]; 
    assign out[4417] = layer_0[3433] ^ layer_0[2270]; 
    assign out[4418] = ~(layer_0[3368] ^ layer_0[7195]); 
    assign out[4419] = ~(layer_0[4770] ^ layer_0[7242]); 
    assign out[4420] = layer_0[1575] ^ layer_0[3266]; 
    assign out[4421] = ~(layer_0[6946] ^ layer_0[7141]); 
    assign out[4422] = ~(layer_0[7874] & layer_0[3487]); 
    assign out[4423] = layer_0[3338]; 
    assign out[4424] = layer_0[104] ^ layer_0[6751]; 
    assign out[4425] = layer_0[6633] ^ layer_0[1747]; 
    assign out[4426] = ~layer_0[2007] | (layer_0[5994] & layer_0[2007]); 
    assign out[4427] = ~(layer_0[7790] ^ layer_0[20]); 
    assign out[4428] = layer_0[146]; 
    assign out[4429] = ~(layer_0[1118] ^ layer_0[7930]); 
    assign out[4430] = layer_0[212]; 
    assign out[4431] = layer_0[1016] ^ layer_0[4280]; 
    assign out[4432] = ~layer_0[6790]; 
    assign out[4433] = ~(layer_0[4423] ^ layer_0[6767]); 
    assign out[4434] = ~layer_0[6992] | (layer_0[4302] & layer_0[6992]); 
    assign out[4435] = layer_0[4188] ^ layer_0[2231]; 
    assign out[4436] = ~layer_0[5993] | (layer_0[107] & layer_0[5993]); 
    assign out[4437] = ~(layer_0[2954] ^ layer_0[6532]); 
    assign out[4438] = ~(layer_0[6687] ^ layer_0[7398]); 
    assign out[4439] = layer_0[562]; 
    assign out[4440] = ~layer_0[3023]; 
    assign out[4441] = ~(layer_0[3609] ^ layer_0[616]); 
    assign out[4442] = layer_0[712] & layer_0[3438]; 
    assign out[4443] = layer_0[7121] | layer_0[3670]; 
    assign out[4444] = ~layer_0[4960] | (layer_0[4960] & layer_0[3857]); 
    assign out[4445] = ~(layer_0[6248] | layer_0[4408]); 
    assign out[4446] = ~layer_0[369] | (layer_0[7506] & layer_0[369]); 
    assign out[4447] = ~layer_0[2865] | (layer_0[2865] & layer_0[3222]); 
    assign out[4448] = ~layer_0[6543] | (layer_0[6543] & layer_0[1809]); 
    assign out[4449] = 1'b1; 
    assign out[4450] = layer_0[1905] | layer_0[2887]; 
    assign out[4451] = ~layer_0[6365]; 
    assign out[4452] = layer_0[4055] ^ layer_0[4124]; 
    assign out[4453] = ~(layer_0[5730] ^ layer_0[7994]); 
    assign out[4454] = ~(layer_0[2943] ^ layer_0[3988]); 
    assign out[4455] = ~(layer_0[1786] ^ layer_0[1977]); 
    assign out[4456] = ~(layer_0[2559] ^ layer_0[4114]); 
    assign out[4457] = ~layer_0[3017] | (layer_0[3017] & layer_0[7647]); 
    assign out[4458] = ~layer_0[4229] | (layer_0[846] & layer_0[4229]); 
    assign out[4459] = ~(layer_0[6113] & layer_0[5705]); 
    assign out[4460] = layer_0[2018]; 
    assign out[4461] = ~(layer_0[1403] & layer_0[2498]); 
    assign out[4462] = ~layer_0[178] | (layer_0[178] & layer_0[1008]); 
    assign out[4463] = ~(layer_0[6015] ^ layer_0[7687]); 
    assign out[4464] = ~(layer_0[4343] & layer_0[3311]); 
    assign out[4465] = ~layer_0[1613] | (layer_0[1613] & layer_0[4147]); 
    assign out[4466] = layer_0[2484] ^ layer_0[3908]; 
    assign out[4467] = ~layer_0[7854]; 
    assign out[4468] = ~layer_0[947]; 
    assign out[4469] = ~layer_0[6387]; 
    assign out[4470] = ~layer_0[1748]; 
    assign out[4471] = layer_0[6488]; 
    assign out[4472] = ~(layer_0[6727] ^ layer_0[990]); 
    assign out[4473] = layer_0[2469] ^ layer_0[2111]; 
    assign out[4474] = layer_0[1749] ^ layer_0[1895]; 
    assign out[4475] = layer_0[481] ^ layer_0[2386]; 
    assign out[4476] = ~layer_0[7618]; 
    assign out[4477] = ~layer_0[759]; 
    assign out[4478] = layer_0[7030]; 
    assign out[4479] = layer_0[4709] ^ layer_0[1615]; 
    assign out[4480] = ~layer_0[1810] | (layer_0[1810] & layer_0[26]); 
    assign out[4481] = layer_0[1131]; 
    assign out[4482] = ~(layer_0[4733] ^ layer_0[6740]); 
    assign out[4483] = ~layer_0[2289]; 
    assign out[4484] = ~layer_0[3189]; 
    assign out[4485] = ~(layer_0[1768] ^ layer_0[5991]); 
    assign out[4486] = ~layer_0[6677] | (layer_0[7494] & layer_0[6677]); 
    assign out[4487] = layer_0[3535] ^ layer_0[2201]; 
    assign out[4488] = layer_0[5190] ^ layer_0[1858]; 
    assign out[4489] = layer_0[347] ^ layer_0[2280]; 
    assign out[4490] = layer_0[3396] ^ layer_0[6957]; 
    assign out[4491] = ~layer_0[4626]; 
    assign out[4492] = layer_0[4394] ^ layer_0[5854]; 
    assign out[4493] = layer_0[3051] & ~layer_0[3663]; 
    assign out[4494] = ~layer_0[6030]; 
    assign out[4495] = layer_0[7722] ^ layer_0[5695]; 
    assign out[4496] = layer_0[4392] | layer_0[3801]; 
    assign out[4497] = layer_0[3006] & layer_0[4303]; 
    assign out[4498] = layer_0[7739] ^ layer_0[1504]; 
    assign out[4499] = ~(layer_0[5889] ^ layer_0[6990]); 
    assign out[4500] = layer_0[5242]; 
    assign out[4501] = layer_0[3058]; 
    assign out[4502] = ~(layer_0[885] ^ layer_0[2470]); 
    assign out[4503] = ~(layer_0[5001] & layer_0[1736]); 
    assign out[4504] = ~layer_0[3950]; 
    assign out[4505] = ~(layer_0[3168] ^ layer_0[2677]); 
    assign out[4506] = ~layer_0[2575]; 
    assign out[4507] = ~(layer_0[4475] ^ layer_0[4981]); 
    assign out[4508] = layer_0[7381] ^ layer_0[5216]; 
    assign out[4509] = ~(layer_0[7919] ^ layer_0[2401]); 
    assign out[4510] = ~(layer_0[10] ^ layer_0[1751]); 
    assign out[4511] = ~(layer_0[3919] ^ layer_0[3825]); 
    assign out[4512] = ~layer_0[1733] | (layer_0[4745] & layer_0[1733]); 
    assign out[4513] = ~layer_0[6108]; 
    assign out[4514] = ~layer_0[2552] | (layer_0[2552] & layer_0[5481]); 
    assign out[4515] = layer_0[3406] ^ layer_0[6585]; 
    assign out[4516] = layer_0[2867] | layer_0[5888]; 
    assign out[4517] = layer_0[7884] ^ layer_0[1938]; 
    assign out[4518] = layer_0[3282]; 
    assign out[4519] = layer_0[1196] ^ layer_0[2943]; 
    assign out[4520] = layer_0[5992] ^ layer_0[7952]; 
    assign out[4521] = layer_0[7218] ^ layer_0[4717]; 
    assign out[4522] = layer_0[1847] ^ layer_0[7762]; 
    assign out[4523] = layer_0[3756]; 
    assign out[4524] = ~(layer_0[7049] ^ layer_0[5608]); 
    assign out[4525] = ~(layer_0[2420] ^ layer_0[7293]); 
    assign out[4526] = ~(layer_0[7822] ^ layer_0[4806]); 
    assign out[4527] = layer_0[5891] ^ layer_0[127]; 
    assign out[4528] = layer_0[307] ^ layer_0[5007]; 
    assign out[4529] = ~layer_0[984] | (layer_0[984] & layer_0[7785]); 
    assign out[4530] = layer_0[6461] ^ layer_0[6139]; 
    assign out[4531] = ~(layer_0[2906] | layer_0[6389]); 
    assign out[4532] = layer_0[3598] ^ layer_0[5198]; 
    assign out[4533] = ~(layer_0[3796] ^ layer_0[7696]); 
    assign out[4534] = ~(layer_0[1814] ^ layer_0[2697]); 
    assign out[4535] = layer_0[7531]; 
    assign out[4536] = ~layer_0[2485]; 
    assign out[4537] = ~(layer_0[3696] & layer_0[3654]); 
    assign out[4538] = ~(layer_0[7643] ^ layer_0[1594]); 
    assign out[4539] = layer_0[7474] & layer_0[5270]; 
    assign out[4540] = ~(layer_0[2221] ^ layer_0[5750]); 
    assign out[4541] = ~layer_0[3536] | (layer_0[3536] & layer_0[3061]); 
    assign out[4542] = layer_0[7512] ^ layer_0[6574]; 
    assign out[4543] = ~layer_0[3251] | (layer_0[3251] & layer_0[1721]); 
    assign out[4544] = layer_0[2327]; 
    assign out[4545] = layer_0[859] | layer_0[5304]; 
    assign out[4546] = layer_0[5417] | layer_0[159]; 
    assign out[4547] = layer_0[4142] & layer_0[2747]; 
    assign out[4548] = layer_0[5003]; 
    assign out[4549] = ~(layer_0[246] ^ layer_0[1780]); 
    assign out[4550] = ~(layer_0[255] ^ layer_0[199]); 
    assign out[4551] = ~(layer_0[3914] & layer_0[2061]); 
    assign out[4552] = layer_0[5542] ^ layer_0[1559]; 
    assign out[4553] = layer_0[2782]; 
    assign out[4554] = layer_0[211] ^ layer_0[3106]; 
    assign out[4555] = ~layer_0[5278]; 
    assign out[4556] = ~layer_0[2824]; 
    assign out[4557] = layer_0[1880] | layer_0[3485]; 
    assign out[4558] = layer_0[2361] & ~layer_0[3130]; 
    assign out[4559] = ~layer_0[5291]; 
    assign out[4560] = layer_0[2369] ^ layer_0[3098]; 
    assign out[4561] = layer_0[7650]; 
    assign out[4562] = ~(layer_0[4610] | layer_0[376]); 
    assign out[4563] = ~(layer_0[5836] ^ layer_0[2692]); 
    assign out[4564] = layer_0[2314] | layer_0[2649]; 
    assign out[4565] = ~(layer_0[7598] & layer_0[6600]); 
    assign out[4566] = layer_0[5657] ^ layer_0[5266]; 
    assign out[4567] = layer_0[82] & ~layer_0[7773]; 
    assign out[4568] = ~(layer_0[2415] ^ layer_0[2426]); 
    assign out[4569] = layer_0[5912] ^ layer_0[6356]; 
    assign out[4570] = layer_0[7964] ^ layer_0[3913]; 
    assign out[4571] = ~(layer_0[3231] & layer_0[33]); 
    assign out[4572] = ~layer_0[128]; 
    assign out[4573] = ~(layer_0[892] & layer_0[6644]); 
    assign out[4574] = ~(layer_0[3458] | layer_0[6208]); 
    assign out[4575] = ~(layer_0[30] ^ layer_0[1917]); 
    assign out[4576] = ~(layer_0[1201] ^ layer_0[1211]); 
    assign out[4577] = ~(layer_0[1079] ^ layer_0[4069]); 
    assign out[4578] = layer_0[3340]; 
    assign out[4579] = ~layer_0[5615] | (layer_0[6690] & layer_0[5615]); 
    assign out[4580] = ~layer_0[2188] | (layer_0[2188] & layer_0[4895]); 
    assign out[4581] = ~(layer_0[6385] ^ layer_0[1903]); 
    assign out[4582] = ~(layer_0[4333] & layer_0[5076]); 
    assign out[4583] = ~(layer_0[3969] ^ layer_0[5540]); 
    assign out[4584] = layer_0[5917] & ~layer_0[691]; 
    assign out[4585] = ~layer_0[2117]; 
    assign out[4586] = ~layer_0[565]; 
    assign out[4587] = ~layer_0[4773]; 
    assign out[4588] = ~(layer_0[918] & layer_0[3252]); 
    assign out[4589] = layer_0[1717]; 
    assign out[4590] = layer_0[3312] | layer_0[451]; 
    assign out[4591] = layer_0[5379] | layer_0[2089]; 
    assign out[4592] = ~(layer_0[7999] ^ layer_0[580]); 
    assign out[4593] = ~layer_0[4045]; 
    assign out[4594] = layer_0[3679] ^ layer_0[6463]; 
    assign out[4595] = ~(layer_0[7582] ^ layer_0[5817]); 
    assign out[4596] = layer_0[6060] ^ layer_0[4124]; 
    assign out[4597] = ~(layer_0[1836] ^ layer_0[6289]); 
    assign out[4598] = layer_0[3026] ^ layer_0[511]; 
    assign out[4599] = layer_0[7626] ^ layer_0[4293]; 
    assign out[4600] = ~layer_0[2153] | (layer_0[1424] & layer_0[2153]); 
    assign out[4601] = ~(layer_0[384] ^ layer_0[5531]); 
    assign out[4602] = layer_0[1693] & ~layer_0[6117]; 
    assign out[4603] = layer_0[2290] & ~layer_0[1193]; 
    assign out[4604] = layer_0[888] & layer_0[7819]; 
    assign out[4605] = ~layer_0[4150] | (layer_0[17] & layer_0[4150]); 
    assign out[4606] = layer_0[6930]; 
    assign out[4607] = ~layer_0[3517] | (layer_0[6777] & layer_0[3517]); 
    assign out[4608] = ~layer_0[6063] | (layer_0[1485] & layer_0[6063]); 
    assign out[4609] = ~layer_0[7887]; 
    assign out[4610] = layer_0[7490] & ~layer_0[3095]; 
    assign out[4611] = layer_0[2104] & ~layer_0[2451]; 
    assign out[4612] = layer_0[2355] ^ layer_0[4482]; 
    assign out[4613] = layer_0[793] ^ layer_0[6847]; 
    assign out[4614] = ~layer_0[7726]; 
    assign out[4615] = ~layer_0[7164] | (layer_0[7164] & layer_0[1146]); 
    assign out[4616] = layer_0[2776] & layer_0[3901]; 
    assign out[4617] = ~(layer_0[6837] ^ layer_0[6014]); 
    assign out[4618] = layer_0[3712] & ~layer_0[7518]; 
    assign out[4619] = layer_0[1624]; 
    assign out[4620] = layer_0[3042] | layer_0[50]; 
    assign out[4621] = layer_0[1620]; 
    assign out[4622] = layer_0[7247] | layer_0[5393]; 
    assign out[4623] = ~(layer_0[5112] ^ layer_0[2787]); 
    assign out[4624] = layer_0[5505] & layer_0[892]; 
    assign out[4625] = ~layer_0[5732]; 
    assign out[4626] = layer_0[3786] & ~layer_0[7022]; 
    assign out[4627] = ~layer_0[5948]; 
    assign out[4628] = layer_0[3271]; 
    assign out[4629] = layer_0[5396] & layer_0[768]; 
    assign out[4630] = layer_0[1526] ^ layer_0[2983]; 
    assign out[4631] = layer_0[3693] & ~layer_0[4244]; 
    assign out[4632] = layer_0[6660] & ~layer_0[4418]; 
    assign out[4633] = layer_0[3562]; 
    assign out[4634] = ~(layer_0[4207] ^ layer_0[1898]); 
    assign out[4635] = layer_0[5914] & layer_0[1581]; 
    assign out[4636] = ~(layer_0[2924] ^ layer_0[5098]); 
    assign out[4637] = layer_0[5533] ^ layer_0[7180]; 
    assign out[4638] = layer_0[4319] & ~layer_0[6364]; 
    assign out[4639] = layer_0[2166] & layer_0[2110]; 
    assign out[4640] = ~layer_0[1546]; 
    assign out[4641] = layer_0[7972] & ~layer_0[2866]; 
    assign out[4642] = ~layer_0[7501] | (layer_0[5155] & layer_0[7501]); 
    assign out[4643] = layer_0[2097] ^ layer_0[5643]; 
    assign out[4644] = layer_0[3891] | layer_0[4441]; 
    assign out[4645] = layer_0[3332] ^ layer_0[4051]; 
    assign out[4646] = ~(layer_0[1090] | layer_0[6206]); 
    assign out[4647] = ~(layer_0[7105] | layer_0[7317]); 
    assign out[4648] = ~(layer_0[1320] & layer_0[7943]); 
    assign out[4649] = ~(layer_0[4485] ^ layer_0[5033]); 
    assign out[4650] = layer_0[5969]; 
    assign out[4651] = ~layer_0[6994]; 
    assign out[4652] = ~(layer_0[7285] | layer_0[7926]); 
    assign out[4653] = layer_0[7598] & ~layer_0[3495]; 
    assign out[4654] = ~(layer_0[2411] ^ layer_0[7088]); 
    assign out[4655] = layer_0[4291] | layer_0[482]; 
    assign out[4656] = ~layer_0[494]; 
    assign out[4657] = ~(layer_0[175] ^ layer_0[5950]); 
    assign out[4658] = layer_0[2107] & ~layer_0[6702]; 
    assign out[4659] = layer_0[2751] ^ layer_0[2432]; 
    assign out[4660] = layer_0[4286] & layer_0[6733]; 
    assign out[4661] = layer_0[5776] & layer_0[4932]; 
    assign out[4662] = layer_0[7356] & ~layer_0[601]; 
    assign out[4663] = ~(layer_0[2127] | layer_0[6341]); 
    assign out[4664] = layer_0[3360] | layer_0[2609]; 
    assign out[4665] = layer_0[5569] & layer_0[3713]; 
    assign out[4666] = layer_0[4504] | layer_0[459]; 
    assign out[4667] = ~(layer_0[7932] ^ layer_0[311]); 
    assign out[4668] = layer_0[89] ^ layer_0[4666]; 
    assign out[4669] = layer_0[4788] ^ layer_0[1574]; 
    assign out[4670] = layer_0[3364] & ~layer_0[1987]; 
    assign out[4671] = ~(layer_0[3941] ^ layer_0[6980]); 
    assign out[4672] = layer_0[1228] & ~layer_0[3979]; 
    assign out[4673] = ~(layer_0[3359] ^ layer_0[1801]); 
    assign out[4674] = ~(layer_0[7220] | layer_0[3103]); 
    assign out[4675] = layer_0[1783] & ~layer_0[5368]; 
    assign out[4676] = ~layer_0[4424] | (layer_0[4424] & layer_0[6698]); 
    assign out[4677] = ~(layer_0[1733] | layer_0[7374]); 
    assign out[4678] = ~layer_0[6741]; 
    assign out[4679] = layer_0[5626] ^ layer_0[7830]; 
    assign out[4680] = layer_0[3447] & layer_0[4506]; 
    assign out[4681] = ~layer_0[5614]; 
    assign out[4682] = ~layer_0[932]; 
    assign out[4683] = ~(layer_0[1886] ^ layer_0[2435]); 
    assign out[4684] = ~(layer_0[5195] | layer_0[3128]); 
    assign out[4685] = layer_0[5013] ^ layer_0[6637]; 
    assign out[4686] = layer_0[2324] ^ layer_0[1645]; 
    assign out[4687] = layer_0[7581]; 
    assign out[4688] = ~layer_0[2884]; 
    assign out[4689] = layer_0[2914]; 
    assign out[4690] = ~(layer_0[6872] ^ layer_0[7677]); 
    assign out[4691] = layer_0[5433]; 
    assign out[4692] = layer_0[7252] & ~layer_0[4865]; 
    assign out[4693] = ~(layer_0[7099] & layer_0[6538]); 
    assign out[4694] = ~(layer_0[2929] ^ layer_0[5629]); 
    assign out[4695] = layer_0[96] | layer_0[6680]; 
    assign out[4696] = layer_0[2994]; 
    assign out[4697] = layer_0[7465] & layer_0[5931]; 
    assign out[4698] = ~layer_0[4184] | (layer_0[2521] & layer_0[4184]); 
    assign out[4699] = ~(layer_0[5894] | layer_0[4326]); 
    assign out[4700] = ~layer_0[7679]; 
    assign out[4701] = ~(layer_0[5922] ^ layer_0[7960]); 
    assign out[4702] = ~(layer_0[5960] ^ layer_0[2656]); 
    assign out[4703] = layer_0[4907] & ~layer_0[4347]; 
    assign out[4704] = layer_0[5617]; 
    assign out[4705] = ~layer_0[4074]; 
    assign out[4706] = ~(layer_0[922] ^ layer_0[3243]); 
    assign out[4707] = layer_0[4902]; 
    assign out[4708] = ~layer_0[7418] | (layer_0[7418] & layer_0[5220]); 
    assign out[4709] = layer_0[7239] ^ layer_0[5804]; 
    assign out[4710] = layer_0[5455] & ~layer_0[6801]; 
    assign out[4711] = ~(layer_0[6089] ^ layer_0[5165]); 
    assign out[4712] = ~(layer_0[2461] ^ layer_0[4720]); 
    assign out[4713] = ~layer_0[5362]; 
    assign out[4714] = layer_0[7619] & ~layer_0[2279]; 
    assign out[4715] = ~(layer_0[3208] ^ layer_0[716]); 
    assign out[4716] = ~(layer_0[5665] | layer_0[5224]); 
    assign out[4717] = ~(layer_0[80] | layer_0[1078]); 
    assign out[4718] = layer_0[2988] & ~layer_0[2357]; 
    assign out[4719] = ~layer_0[5672]; 
    assign out[4720] = layer_0[7201] ^ layer_0[7924]; 
    assign out[4721] = ~(layer_0[2527] | layer_0[4578]); 
    assign out[4722] = ~(layer_0[4893] | layer_0[5074]); 
    assign out[4723] = layer_0[1678]; 
    assign out[4724] = ~layer_0[3164]; 
    assign out[4725] = ~(layer_0[5648] & layer_0[5739]); 
    assign out[4726] = ~(layer_0[1752] ^ layer_0[3893]); 
    assign out[4727] = ~(layer_0[2689] ^ layer_0[6705]); 
    assign out[4728] = layer_0[833] & ~layer_0[53]; 
    assign out[4729] = layer_0[1166] ^ layer_0[3383]; 
    assign out[4730] = ~(layer_0[5093] ^ layer_0[4646]); 
    assign out[4731] = layer_0[1291]; 
    assign out[4732] = layer_0[5374] & layer_0[6417]; 
    assign out[4733] = layer_0[3759] & ~layer_0[7585]; 
    assign out[4734] = ~layer_0[5731]; 
    assign out[4735] = layer_0[2019] & layer_0[1820]; 
    assign out[4736] = layer_0[2510] ^ layer_0[1433]; 
    assign out[4737] = layer_0[5815] & ~layer_0[2025]; 
    assign out[4738] = ~layer_0[3021]; 
    assign out[4739] = ~layer_0[2712]; 
    assign out[4740] = ~layer_0[595] | (layer_0[595] & layer_0[2792]); 
    assign out[4741] = layer_0[2997] | layer_0[1767]; 
    assign out[4742] = layer_0[5808] ^ layer_0[6135]; 
    assign out[4743] = ~(layer_0[3109] ^ layer_0[729]); 
    assign out[4744] = ~layer_0[4359]; 
    assign out[4745] = layer_0[7556] ^ layer_0[4628]; 
    assign out[4746] = ~layer_0[2022]; 
    assign out[4747] = layer_0[883] & ~layer_0[1611]; 
    assign out[4748] = layer_0[6564] & ~layer_0[7826]; 
    assign out[4749] = layer_0[3382] & ~layer_0[2408]; 
    assign out[4750] = layer_0[5693]; 
    assign out[4751] = layer_0[1663]; 
    assign out[4752] = layer_0[7877] & ~layer_0[7475]; 
    assign out[4753] = layer_0[470]; 
    assign out[4754] = layer_0[1241] & layer_0[2968]; 
    assign out[4755] = ~(layer_0[3427] ^ layer_0[2307]); 
    assign out[4756] = ~layer_0[1704]; 
    assign out[4757] = layer_0[3563] & ~layer_0[855]; 
    assign out[4758] = ~(layer_0[1466] ^ layer_0[2270]); 
    assign out[4759] = ~(layer_0[392] | layer_0[873]); 
    assign out[4760] = ~layer_0[2623]; 
    assign out[4761] = ~(layer_0[5179] ^ layer_0[3136]); 
    assign out[4762] = ~(layer_0[1090] | layer_0[7683]); 
    assign out[4763] = ~layer_0[6392] | (layer_0[6392] & layer_0[5504]); 
    assign out[4764] = layer_0[7843] & ~layer_0[6372]; 
    assign out[4765] = ~(layer_0[6456] ^ layer_0[7536]); 
    assign out[4766] = layer_0[3063]; 
    assign out[4767] = layer_0[6350] & layer_0[2661]; 
    assign out[4768] = ~(layer_0[6184] ^ layer_0[1462]); 
    assign out[4769] = ~(layer_0[4412] | layer_0[7709]); 
    assign out[4770] = ~(layer_0[927] | layer_0[2410]); 
    assign out[4771] = layer_0[7513] & layer_0[4235]; 
    assign out[4772] = ~(layer_0[1363] ^ layer_0[1428]); 
    assign out[4773] = layer_0[956]; 
    assign out[4774] = layer_0[4063] & ~layer_0[4353]; 
    assign out[4775] = layer_0[5737] & ~layer_0[150]; 
    assign out[4776] = ~(layer_0[5068] | layer_0[4183]); 
    assign out[4777] = ~layer_0[7340] | (layer_0[493] & layer_0[7340]); 
    assign out[4778] = layer_0[7810] & ~layer_0[6247]; 
    assign out[4779] = layer_0[2613] ^ layer_0[3169]; 
    assign out[4780] = layer_0[85] & layer_0[6019]; 
    assign out[4781] = layer_0[2129] & ~layer_0[636]; 
    assign out[4782] = layer_0[5569] & layer_0[2549]; 
    assign out[4783] = layer_0[7602] & ~layer_0[6422]; 
    assign out[4784] = ~(layer_0[4222] ^ layer_0[560]); 
    assign out[4785] = ~layer_0[2724] | (layer_0[5201] & layer_0[2724]); 
    assign out[4786] = ~layer_0[2090] | (layer_0[3974] & layer_0[2090]); 
    assign out[4787] = layer_0[2262] ^ layer_0[1110]; 
    assign out[4788] = layer_0[3379] ^ layer_0[5245]; 
    assign out[4789] = layer_0[6358] ^ layer_0[7876]; 
    assign out[4790] = layer_0[198] & layer_0[7439]; 
    assign out[4791] = ~(layer_0[6283] ^ layer_0[695]); 
    assign out[4792] = layer_0[5265]; 
    assign out[4793] = ~(layer_0[5144] ^ layer_0[5230]); 
    assign out[4794] = layer_0[2039] & ~layer_0[230]; 
    assign out[4795] = ~(layer_0[3529] ^ layer_0[2167]); 
    assign out[4796] = ~(layer_0[661] | layer_0[3136]); 
    assign out[4797] = layer_0[416] & ~layer_0[1014]; 
    assign out[4798] = layer_0[358]; 
    assign out[4799] = ~layer_0[4227]; 
    assign out[4800] = ~(layer_0[4941] & layer_0[6759]); 
    assign out[4801] = layer_0[2563] ^ layer_0[2874]; 
    assign out[4802] = layer_0[5500] & layer_0[5843]; 
    assign out[4803] = ~(layer_0[4043] ^ layer_0[5594]); 
    assign out[4804] = ~(layer_0[4438] ^ layer_0[220]); 
    assign out[4805] = ~layer_0[5968]; 
    assign out[4806] = ~(layer_0[4091] ^ layer_0[2713]); 
    assign out[4807] = layer_0[1063]; 
    assign out[4808] = ~(layer_0[4107] & layer_0[3950]); 
    assign out[4809] = ~layer_0[7631]; 
    assign out[4810] = layer_0[5174] & layer_0[7212]; 
    assign out[4811] = layer_0[1395] & layer_0[5734]; 
    assign out[4812] = layer_0[5604]; 
    assign out[4813] = layer_0[889]; 
    assign out[4814] = layer_0[6736]; 
    assign out[4815] = layer_0[2820] & layer_0[2944]; 
    assign out[4816] = layer_0[3179]; 
    assign out[4817] = layer_0[6880] ^ layer_0[1800]; 
    assign out[4818] = layer_0[1906]; 
    assign out[4819] = ~(layer_0[7863] & layer_0[7261]); 
    assign out[4820] = layer_0[2561]; 
    assign out[4821] = layer_0[7451]; 
    assign out[4822] = ~(layer_0[5256] | layer_0[6805]); 
    assign out[4823] = ~(layer_0[5285] ^ layer_0[618]); 
    assign out[4824] = ~(layer_0[6716] | layer_0[1747]); 
    assign out[4825] = ~(layer_0[2136] ^ layer_0[6091]); 
    assign out[4826] = layer_0[2] | layer_0[3858]; 
    assign out[4827] = ~(layer_0[5925] ^ layer_0[3171]); 
    assign out[4828] = ~layer_0[3303]; 
    assign out[4829] = layer_0[1690] & layer_0[7263]; 
    assign out[4830] = layer_0[7230] ^ layer_0[7711]; 
    assign out[4831] = layer_0[4538] ^ layer_0[1520]; 
    assign out[4832] = layer_0[7357] ^ layer_0[3975]; 
    assign out[4833] = ~(layer_0[2087] ^ layer_0[2420]); 
    assign out[4834] = ~(layer_0[1490] ^ layer_0[3422]); 
    assign out[4835] = layer_0[7956] & layer_0[5432]; 
    assign out[4836] = ~layer_0[58]; 
    assign out[4837] = layer_0[5412] ^ layer_0[3916]; 
    assign out[4838] = layer_0[5787] & layer_0[4175]; 
    assign out[4839] = layer_0[4785]; 
    assign out[4840] = layer_0[6163] | layer_0[5511]; 
    assign out[4841] = ~layer_0[2569]; 
    assign out[4842] = layer_0[3177] ^ layer_0[2338]; 
    assign out[4843] = layer_0[153]; 
    assign out[4844] = ~layer_0[713]; 
    assign out[4845] = ~(layer_0[5628] | layer_0[6176]); 
    assign out[4846] = layer_0[1932] & layer_0[2146]; 
    assign out[4847] = layer_0[7699]; 
    assign out[4848] = layer_0[567] & ~layer_0[4275]; 
    assign out[4849] = layer_0[4715] & ~layer_0[1337]; 
    assign out[4850] = ~layer_0[5859]; 
    assign out[4851] = layer_0[867]; 
    assign out[4852] = ~(layer_0[2668] ^ layer_0[2002]); 
    assign out[4853] = ~layer_0[2828]; 
    assign out[4854] = ~(layer_0[3478] ^ layer_0[3238]); 
    assign out[4855] = layer_0[5452] & layer_0[5313]; 
    assign out[4856] = layer_0[784] & ~layer_0[656]; 
    assign out[4857] = ~layer_0[7737]; 
    assign out[4858] = layer_0[5751] ^ layer_0[1591]; 
    assign out[4859] = ~(layer_0[7871] | layer_0[2984]); 
    assign out[4860] = ~layer_0[4659]; 
    assign out[4861] = ~layer_0[2308]; 
    assign out[4862] = ~(layer_0[2182] ^ layer_0[2436]); 
    assign out[4863] = ~(layer_0[7653] | layer_0[7031]); 
    assign out[4864] = layer_0[7234] & ~layer_0[7480]; 
    assign out[4865] = layer_0[3119] ^ layer_0[2663]; 
    assign out[4866] = ~(layer_0[4660] | layer_0[5348]); 
    assign out[4867] = layer_0[7105] | layer_0[791]; 
    assign out[4868] = layer_0[1253] ^ layer_0[6959]; 
    assign out[4869] = layer_0[267] & ~layer_0[6160]; 
    assign out[4870] = layer_0[6989] & layer_0[6494]; 
    assign out[4871] = layer_0[3123] | layer_0[6434]; 
    assign out[4872] = ~(layer_0[2926] ^ layer_0[5554]); 
    assign out[4873] = layer_0[3475] ^ layer_0[6503]; 
    assign out[4874] = layer_0[6603] & ~layer_0[5853]; 
    assign out[4875] = ~layer_0[5715] | (layer_0[1401] & layer_0[5715]); 
    assign out[4876] = layer_0[4887]; 
    assign out[4877] = ~(layer_0[7022] ^ layer_0[7196]); 
    assign out[4878] = ~layer_0[7927] | (layer_0[6363] & layer_0[7927]); 
    assign out[4879] = layer_0[5010] | layer_0[4750]; 
    assign out[4880] = ~layer_0[262]; 
    assign out[4881] = layer_0[2948] ^ layer_0[7534]; 
    assign out[4882] = ~(layer_0[4846] | layer_0[7707]); 
    assign out[4883] = layer_0[2583] ^ layer_0[6344]; 
    assign out[4884] = layer_0[4974] | layer_0[5707]; 
    assign out[4885] = ~(layer_0[5142] ^ layer_0[5255]); 
    assign out[4886] = ~(layer_0[6127] | layer_0[966]); 
    assign out[4887] = ~(layer_0[5773] | layer_0[5369]); 
    assign out[4888] = ~(layer_0[3030] ^ layer_0[740]); 
    assign out[4889] = layer_0[6830] & ~layer_0[256]; 
    assign out[4890] = ~(layer_0[1725] ^ layer_0[3697]); 
    assign out[4891] = layer_0[4935]; 
    assign out[4892] = ~(layer_0[3259] ^ layer_0[1596]); 
    assign out[4893] = layer_0[1278]; 
    assign out[4894] = ~(layer_0[3913] ^ layer_0[6488]); 
    assign out[4895] = layer_0[6246] ^ layer_0[1365]; 
    assign out[4896] = ~(layer_0[577] ^ layer_0[5002]); 
    assign out[4897] = layer_0[3856] & ~layer_0[7192]; 
    assign out[4898] = layer_0[1115] & ~layer_0[7255]; 
    assign out[4899] = layer_0[1958] & layer_0[202]; 
    assign out[4900] = layer_0[6755]; 
    assign out[4901] = ~layer_0[221]; 
    assign out[4902] = layer_0[4982] & layer_0[7735]; 
    assign out[4903] = ~layer_0[6877]; 
    assign out[4904] = ~(layer_0[2848] | layer_0[5424]); 
    assign out[4905] = ~(layer_0[3589] ^ layer_0[7119]); 
    assign out[4906] = layer_0[7102] & ~layer_0[700]; 
    assign out[4907] = layer_0[4729]; 
    assign out[4908] = layer_0[2758] ^ layer_0[6757]; 
    assign out[4909] = layer_0[4784]; 
    assign out[4910] = ~layer_0[2287] | (layer_0[2287] & layer_0[2184]); 
    assign out[4911] = layer_0[387]; 
    assign out[4912] = layer_0[7295] ^ layer_0[580]; 
    assign out[4913] = layer_0[88] ^ layer_0[3184]; 
    assign out[4914] = layer_0[4060] ^ layer_0[4270]; 
    assign out[4915] = layer_0[495] | layer_0[4555]; 
    assign out[4916] = layer_0[5072] ^ layer_0[403]; 
    assign out[4917] = layer_0[4830] ^ layer_0[219]; 
    assign out[4918] = layer_0[4847] & ~layer_0[24]; 
    assign out[4919] = ~(layer_0[5383] & layer_0[1051]); 
    assign out[4920] = layer_0[375] & ~layer_0[6271]; 
    assign out[4921] = ~(layer_0[3554] ^ layer_0[4513]); 
    assign out[4922] = layer_0[5083] & ~layer_0[3166]; 
    assign out[4923] = ~(layer_0[1114] ^ layer_0[1203]); 
    assign out[4924] = ~layer_0[4063]; 
    assign out[4925] = layer_0[5020] | layer_0[7865]; 
    assign out[4926] = layer_0[6974] ^ layer_0[1468]; 
    assign out[4927] = ~(layer_0[6486] ^ layer_0[7589]); 
    assign out[4928] = layer_0[2279] ^ layer_0[6810]; 
    assign out[4929] = ~layer_0[3486]; 
    assign out[4930] = layer_0[413] ^ layer_0[6984]; 
    assign out[4931] = layer_0[4970] ^ layer_0[5828]; 
    assign out[4932] = layer_0[6459] & ~layer_0[7244]; 
    assign out[4933] = ~(layer_0[4829] ^ layer_0[6168]); 
    assign out[4934] = layer_0[7021] | layer_0[707]; 
    assign out[4935] = ~layer_0[734]; 
    assign out[4936] = layer_0[6879] & layer_0[5476]; 
    assign out[4937] = ~layer_0[5171]; 
    assign out[4938] = layer_0[70] & layer_0[5946]; 
    assign out[4939] = ~(layer_0[4532] ^ layer_0[2958]); 
    assign out[4940] = layer_0[1919]; 
    assign out[4941] = ~layer_0[7745] | (layer_0[7882] & layer_0[7745]); 
    assign out[4942] = layer_0[2528]; 
    assign out[4943] = layer_0[2329] ^ layer_0[3955]; 
    assign out[4944] = ~(layer_0[4825] | layer_0[7296]); 
    assign out[4945] = layer_0[6579] ^ layer_0[1339]; 
    assign out[4946] = layer_0[7172] ^ layer_0[2670]; 
    assign out[4947] = layer_0[3301] & layer_0[1666]; 
    assign out[4948] = layer_0[639]; 
    assign out[4949] = layer_0[5658] ^ layer_0[1457]; 
    assign out[4950] = ~layer_0[122]; 
    assign out[4951] = layer_0[1541] ^ layer_0[3604]; 
    assign out[4952] = ~(layer_0[2297] ^ layer_0[3215]); 
    assign out[4953] = layer_0[1288] & ~layer_0[321]; 
    assign out[4954] = ~(layer_0[4188] | layer_0[3203]); 
    assign out[4955] = ~(layer_0[1974] | layer_0[5122]); 
    assign out[4956] = ~layer_0[3552]; 
    assign out[4957] = ~(layer_0[5152] ^ layer_0[2621]); 
    assign out[4958] = layer_0[1790] ^ layer_0[4286]; 
    assign out[4959] = layer_0[7474] & layer_0[7712]; 
    assign out[4960] = layer_0[3002] ^ layer_0[4695]; 
    assign out[4961] = layer_0[1997] & ~layer_0[1320]; 
    assign out[4962] = layer_0[6157] & ~layer_0[166]; 
    assign out[4963] = layer_0[555] & ~layer_0[2196]; 
    assign out[4964] = layer_0[7058]; 
    assign out[4965] = layer_0[5559]; 
    assign out[4966] = layer_0[3186] ^ layer_0[331]; 
    assign out[4967] = layer_0[2048] ^ layer_0[3190]; 
    assign out[4968] = layer_0[269] & ~layer_0[7723]; 
    assign out[4969] = layer_0[2606] | layer_0[954]; 
    assign out[4970] = layer_0[760] & layer_0[7249]; 
    assign out[4971] = ~layer_0[4859] | (layer_0[469] & layer_0[4859]); 
    assign out[4972] = ~(layer_0[7412] ^ layer_0[5329]); 
    assign out[4973] = layer_0[5054] ^ layer_0[5140]; 
    assign out[4974] = layer_0[834] & ~layer_0[6072]; 
    assign out[4975] = layer_0[1484] & ~layer_0[5519]; 
    assign out[4976] = ~layer_0[4480]; 
    assign out[4977] = ~(layer_0[2882] | layer_0[1332]); 
    assign out[4978] = layer_0[7651] ^ layer_0[142]; 
    assign out[4979] = layer_0[5032]; 
    assign out[4980] = ~layer_0[73]; 
    assign out[4981] = layer_0[1297] & layer_0[5862]; 
    assign out[4982] = ~(layer_0[3927] ^ layer_0[6291]); 
    assign out[4983] = layer_0[3848] | layer_0[3267]; 
    assign out[4984] = ~layer_0[5859]; 
    assign out[4985] = layer_0[4026]; 
    assign out[4986] = ~(layer_0[3217] ^ layer_0[6119]); 
    assign out[4987] = ~(layer_0[736] | layer_0[3284]); 
    assign out[4988] = layer_0[4121]; 
    assign out[4989] = layer_0[3947] & layer_0[826]; 
    assign out[4990] = layer_0[1126] ^ layer_0[7394]; 
    assign out[4991] = layer_0[5180] ^ layer_0[3089]; 
    assign out[4992] = layer_0[4142] ^ layer_0[7539]; 
    assign out[4993] = layer_0[1380]; 
    assign out[4994] = ~(layer_0[3646] & layer_0[1599]); 
    assign out[4995] = ~(layer_0[6190] | layer_0[4812]); 
    assign out[4996] = layer_0[2581]; 
    assign out[4997] = layer_0[1634] ^ layer_0[3681]; 
    assign out[4998] = layer_0[2354]; 
    assign out[4999] = layer_0[6570] ^ layer_0[4332]; 
    assign out[5000] = ~layer_0[6377]; 
    assign out[5001] = layer_0[5428] & ~layer_0[1328]; 
    assign out[5002] = layer_0[1154] ^ layer_0[5612]; 
    assign out[5003] = layer_0[2266] & layer_0[2632]; 
    assign out[5004] = layer_0[6253] & layer_0[7787]; 
    assign out[5005] = ~(layer_0[5791] ^ layer_0[1287]); 
    assign out[5006] = layer_0[6131] ^ layer_0[7243]; 
    assign out[5007] = ~(layer_0[1942] ^ layer_0[1877]); 
    assign out[5008] = layer_0[4106] ^ layer_0[3992]; 
    assign out[5009] = ~(layer_0[4508] ^ layer_0[2850]); 
    assign out[5010] = layer_0[1582] ^ layer_0[7910]; 
    assign out[5011] = ~(layer_0[513] ^ layer_0[7034]); 
    assign out[5012] = ~(layer_0[4448] | layer_0[4966]); 
    assign out[5013] = ~(layer_0[870] | layer_0[1190]); 
    assign out[5014] = layer_0[2529] | layer_0[2282]; 
    assign out[5015] = ~(layer_0[52] ^ layer_0[3737]); 
    assign out[5016] = ~(layer_0[3889] ^ layer_0[7656]); 
    assign out[5017] = layer_0[116] & layer_0[6997]; 
    assign out[5018] = layer_0[6674] & layer_0[2116]; 
    assign out[5019] = layer_0[4126]; 
    assign out[5020] = ~(layer_0[6513] ^ layer_0[1578]); 
    assign out[5021] = layer_0[7365] & ~layer_0[2179]; 
    assign out[5022] = ~layer_0[5703]; 
    assign out[5023] = ~layer_0[6351]; 
    assign out[5024] = layer_0[3000] & ~layer_0[5264]; 
    assign out[5025] = layer_0[6740] ^ layer_0[6106]; 
    assign out[5026] = layer_0[7292] & ~layer_0[3129]; 
    assign out[5027] = ~(layer_0[5498] | layer_0[6826]); 
    assign out[5028] = ~(layer_0[5804] ^ layer_0[444]); 
    assign out[5029] = layer_0[3944] ^ layer_0[3446]; 
    assign out[5030] = ~layer_0[6947] | (layer_0[6947] & layer_0[6659]); 
    assign out[5031] = ~(layer_0[5718] | layer_0[2770]); 
    assign out[5032] = layer_0[6094] ^ layer_0[5016]; 
    assign out[5033] = layer_0[6729]; 
    assign out[5034] = layer_0[1758]; 
    assign out[5035] = layer_0[4105] & ~layer_0[1845]; 
    assign out[5036] = ~layer_0[2473]; 
    assign out[5037] = ~(layer_0[2714] ^ layer_0[800]); 
    assign out[5038] = layer_0[1520] ^ layer_0[1363]; 
    assign out[5039] = ~(layer_0[3493] | layer_0[710]); 
    assign out[5040] = layer_0[7849]; 
    assign out[5041] = layer_0[1340] & ~layer_0[3400]; 
    assign out[5042] = layer_0[5402] & ~layer_0[6340]; 
    assign out[5043] = layer_0[2790] | layer_0[7920]; 
    assign out[5044] = layer_0[5928] & ~layer_0[5510]; 
    assign out[5045] = ~layer_0[7625] | (layer_0[409] & layer_0[7625]); 
    assign out[5046] = layer_0[6988] & ~layer_0[2014]; 
    assign out[5047] = layer_0[2537]; 
    assign out[5048] = layer_0[4639] & ~layer_0[147]; 
    assign out[5049] = layer_0[4689] & ~layer_0[3920]; 
    assign out[5050] = ~(layer_0[310] & layer_0[4152]); 
    assign out[5051] = layer_0[7974] & layer_0[2323]; 
    assign out[5052] = ~(layer_0[4653] ^ layer_0[997]); 
    assign out[5053] = layer_0[2120]; 
    assign out[5054] = layer_0[3731] ^ layer_0[7019]; 
    assign out[5055] = ~(layer_0[1374] | layer_0[6521]); 
    assign out[5056] = layer_0[2550] & ~layer_0[7347]; 
    assign out[5057] = layer_0[1893]; 
    assign out[5058] = layer_0[2266]; 
    assign out[5059] = layer_0[2192] & ~layer_0[1431]; 
    assign out[5060] = ~layer_0[6612]; 
    assign out[5061] = ~(layer_0[2121] ^ layer_0[6614]); 
    assign out[5062] = layer_0[2100] ^ layer_0[3613]; 
    assign out[5063] = layer_0[617]; 
    assign out[5064] = ~(layer_0[4990] ^ layer_0[2849]); 
    assign out[5065] = layer_0[309] & layer_0[3661]; 
    assign out[5066] = layer_0[638] & ~layer_0[4624]; 
    assign out[5067] = ~(layer_0[5735] ^ layer_0[5361]); 
    assign out[5068] = layer_0[431] & layer_0[805]; 
    assign out[5069] = ~layer_0[1721]; 
    assign out[5070] = ~layer_0[4550]; 
    assign out[5071] = ~(layer_0[7330] ^ layer_0[3285]); 
    assign out[5072] = layer_0[6651] & layer_0[830]; 
    assign out[5073] = layer_0[7945]; 
    assign out[5074] = layer_0[6352] & ~layer_0[4313]; 
    assign out[5075] = ~(layer_0[2812] | layer_0[1139]); 
    assign out[5076] = layer_0[2657] & layer_0[2202]; 
    assign out[5077] = ~(layer_0[6038] ^ layer_0[4432]); 
    assign out[5078] = layer_0[7939] ^ layer_0[619]; 
    assign out[5079] = ~layer_0[2724]; 
    assign out[5080] = ~layer_0[3518] | (layer_0[3000] & layer_0[3518]); 
    assign out[5081] = layer_0[628]; 
    assign out[5082] = layer_0[7520]; 
    assign out[5083] = ~(layer_0[5366] ^ layer_0[5041]); 
    assign out[5084] = layer_0[1290] | layer_0[3986]; 
    assign out[5085] = layer_0[2620] & layer_0[109]; 
    assign out[5086] = ~layer_0[765]; 
    assign out[5087] = ~(layer_0[2947] & layer_0[1502]); 
    assign out[5088] = ~layer_0[51]; 
    assign out[5089] = ~layer_0[4020] | (layer_0[849] & layer_0[4020]); 
    assign out[5090] = ~layer_0[3964]; 
    assign out[5091] = layer_0[5339] ^ layer_0[6322]; 
    assign out[5092] = ~layer_0[1911]; 
    assign out[5093] = ~(layer_0[7216] | layer_0[1435]); 
    assign out[5094] = layer_0[2654] ^ layer_0[1480]; 
    assign out[5095] = ~layer_0[7280] | (layer_0[7280] & layer_0[6282]); 
    assign out[5096] = ~(layer_0[4000] ^ layer_0[690]); 
    assign out[5097] = layer_0[3187] ^ layer_0[397]; 
    assign out[5098] = layer_0[1817] & ~layer_0[3850]; 
    assign out[5099] = ~layer_0[5936]; 
    assign out[5100] = layer_0[4350] ^ layer_0[2603]; 
    assign out[5101] = layer_0[2198] & ~layer_0[3979]; 
    assign out[5102] = layer_0[6591] & ~layer_0[1069]; 
    assign out[5103] = layer_0[6354] ^ layer_0[611]; 
    assign out[5104] = layer_0[5956] ^ layer_0[3011]; 
    assign out[5105] = layer_0[1494] & ~layer_0[3326]; 
    assign out[5106] = layer_0[7151] & ~layer_0[5369]; 
    assign out[5107] = ~layer_0[6943] | (layer_0[1767] & layer_0[6943]); 
    assign out[5108] = layer_0[3886] & layer_0[4297]; 
    assign out[5109] = layer_0[4165] & ~layer_0[3501]; 
    assign out[5110] = 1'b0; 
    assign out[5111] = 1'b0; 
    assign out[5112] = 1'b0; 
    assign out[5113] = 1'b0; 
    assign out[5114] = 1'b0; 
    assign out[5115] = 1'b0; 
    assign out[5116] = 1'b0; 
    assign out[5117] = 1'b0; 
    assign out[5118] = 1'b0; 
    assign out[5119] = 1'b0; 
    assign out[5120] = 1'b0; 
    assign out[5121] = 1'b0; 
    assign out[5122] = 1'b0; 
    assign out[5123] = 1'b0; 
    assign out[5124] = 1'b0; 
    assign out[5125] = 1'b0; 
    assign out[5126] = 1'b0; 
    assign out[5127] = 1'b0; 
    assign out[5128] = 1'b0; 
    assign out[5129] = 1'b0; 
    assign out[5130] = 1'b0; 
    assign out[5131] = 1'b0; 
    assign out[5132] = 1'b0; 
    assign out[5133] = 1'b0; 
    assign out[5134] = 1'b0; 
    assign out[5135] = 1'b0; 
    assign out[5136] = 1'b0; 
    assign out[5137] = 1'b0; 
    assign out[5138] = 1'b0; 
    assign out[5139] = 1'b0; 
    assign out[5140] = 1'b0; 
    assign out[5141] = 1'b0; 
    assign out[5142] = 1'b0; 
    assign out[5143] = 1'b0; 
    assign out[5144] = 1'b0; 
    assign out[5145] = 1'b0; 
    assign out[5146] = 1'b0; 
    assign out[5147] = 1'b0; 
    assign out[5148] = 1'b0; 
    assign out[5149] = 1'b0; 
    assign out[5150] = 1'b0; 
    assign out[5151] = 1'b0; 
    assign out[5152] = 1'b0; 
    assign out[5153] = 1'b0; 
    assign out[5154] = 1'b0; 
    assign out[5155] = 1'b0; 
    assign out[5156] = 1'b0; 
    assign out[5157] = 1'b0; 
    assign out[5158] = 1'b0; 
    assign out[5159] = 1'b0; 
    assign out[5160] = 1'b0; 
    assign out[5161] = 1'b0; 
    assign out[5162] = 1'b0; 
    assign out[5163] = 1'b0; 
    assign out[5164] = 1'b0; 
    assign out[5165] = 1'b0; 
    assign out[5166] = 1'b0; 
    assign out[5167] = 1'b0; 
    assign out[5168] = 1'b0; 
    assign out[5169] = 1'b0; 
    assign out[5170] = 1'b0; 
    assign out[5171] = 1'b0; 
    assign out[5172] = 1'b0; 
    assign out[5173] = 1'b0; 
    assign out[5174] = 1'b0; 
    assign out[5175] = 1'b0; 
    assign out[5176] = 1'b0; 
    assign out[5177] = 1'b0; 
    assign out[5178] = 1'b0; 
    assign out[5179] = 1'b0; 
    assign out[5180] = 1'b0; 
    assign out[5181] = 1'b0; 
    assign out[5182] = 1'b0; 
    assign out[5183] = 1'b0; 
    assign out[5184] = 1'b0; 
    assign out[5185] = 1'b0; 
    assign out[5186] = 1'b0; 
    assign out[5187] = 1'b0; 
    assign out[5188] = 1'b0; 
    assign out[5189] = 1'b0; 
    assign out[5190] = 1'b0; 
    assign out[5191] = 1'b0; 
    assign out[5192] = 1'b0; 
    assign out[5193] = 1'b0; 
    assign out[5194] = 1'b0; 
    assign out[5195] = 1'b0; 
    assign out[5196] = 1'b0; 
    assign out[5197] = 1'b0; 
    assign out[5198] = 1'b0; 
    assign out[5199] = 1'b0; 
    assign out[5200] = 1'b0; 
    assign out[5201] = 1'b0; 
    assign out[5202] = 1'b0; 
    assign out[5203] = 1'b0; 
    assign out[5204] = 1'b0; 
    assign out[5205] = 1'b0; 
    assign out[5206] = 1'b0; 
    assign out[5207] = 1'b0; 
    assign out[5208] = 1'b0; 
    assign out[5209] = 1'b0; 
    assign out[5210] = 1'b0; 
    assign out[5211] = 1'b0; 
    assign out[5212] = 1'b0; 
    assign out[5213] = 1'b0; 
    assign out[5214] = 1'b0; 
    assign out[5215] = 1'b0; 
    assign out[5216] = 1'b0; 
    assign out[5217] = 1'b0; 
    assign out[5218] = 1'b0; 
    assign out[5219] = 1'b0; 
    assign out[5220] = 1'b0; 
    assign out[5221] = 1'b0; 
    assign out[5222] = 1'b0; 
    assign out[5223] = 1'b0; 
    assign out[5224] = 1'b0; 
    assign out[5225] = 1'b0; 
    assign out[5226] = 1'b0; 
    assign out[5227] = 1'b0; 
    assign out[5228] = 1'b0; 
    assign out[5229] = 1'b0; 
    assign out[5230] = 1'b0; 
    assign out[5231] = 1'b0; 
    assign out[5232] = 1'b0; 
    assign out[5233] = 1'b0; 
    assign out[5234] = 1'b0; 
    assign out[5235] = 1'b0; 
    assign out[5236] = 1'b0; 
    assign out[5237] = 1'b0; 
    assign out[5238] = 1'b0; 
    assign out[5239] = 1'b0; 
    assign out[5240] = 1'b0; 
    assign out[5241] = 1'b0; 
    assign out[5242] = 1'b0; 
    assign out[5243] = 1'b0; 
    assign out[5244] = 1'b0; 
    assign out[5245] = 1'b0; 
    assign out[5246] = 1'b0; 
    assign out[5247] = 1'b0; 
    assign out[5248] = 1'b0; 
    assign out[5249] = 1'b0; 
    assign out[5250] = 1'b0; 
    assign out[5251] = 1'b0; 
    assign out[5252] = 1'b0; 
    assign out[5253] = 1'b0; 
    assign out[5254] = 1'b0; 
    assign out[5255] = 1'b0; 
    assign out[5256] = 1'b0; 
    assign out[5257] = 1'b0; 
    assign out[5258] = 1'b0; 
    assign out[5259] = 1'b0; 
    assign out[5260] = 1'b0; 
    assign out[5261] = 1'b0; 
    assign out[5262] = 1'b0; 
    assign out[5263] = 1'b0; 
    assign out[5264] = 1'b0; 
    assign out[5265] = 1'b0; 
    assign out[5266] = 1'b0; 
    assign out[5267] = 1'b0; 
    assign out[5268] = 1'b0; 
    assign out[5269] = 1'b0; 
    assign out[5270] = 1'b0; 
    assign out[5271] = 1'b0; 
    assign out[5272] = 1'b0; 
    assign out[5273] = 1'b0; 
    assign out[5274] = 1'b0; 
    assign out[5275] = 1'b0; 
    assign out[5276] = 1'b0; 
    assign out[5277] = 1'b0; 
    assign out[5278] = 1'b0; 
    assign out[5279] = 1'b0; 
    assign out[5280] = 1'b0; 
    assign out[5281] = 1'b0; 
    assign out[5282] = 1'b0; 
    assign out[5283] = 1'b0; 
    assign out[5284] = 1'b0; 
    assign out[5285] = 1'b0; 
    assign out[5286] = 1'b0; 
    assign out[5287] = 1'b0; 
    assign out[5288] = 1'b0; 
    assign out[5289] = 1'b0; 
    assign out[5290] = 1'b0; 
    assign out[5291] = 1'b0; 
    assign out[5292] = 1'b0; 
    assign out[5293] = 1'b0; 
    assign out[5294] = 1'b0; 
    assign out[5295] = 1'b0; 
    assign out[5296] = 1'b0; 
    assign out[5297] = 1'b0; 
    assign out[5298] = 1'b0; 
    assign out[5299] = 1'b0; 
    assign out[5300] = 1'b0; 
    assign out[5301] = 1'b0; 
    assign out[5302] = 1'b0; 
    assign out[5303] = 1'b0; 
    assign out[5304] = 1'b0; 
    assign out[5305] = 1'b0; 
    assign out[5306] = 1'b0; 
    assign out[5307] = 1'b0; 
    assign out[5308] = 1'b0; 
    assign out[5309] = 1'b0; 
    assign out[5310] = 1'b0; 
    assign out[5311] = 1'b0; 
    assign out[5312] = 1'b0; 
    assign out[5313] = 1'b0; 
    assign out[5314] = 1'b0; 
    assign out[5315] = 1'b0; 
    assign out[5316] = 1'b0; 
    assign out[5317] = 1'b0; 
    assign out[5318] = 1'b0; 
    assign out[5319] = 1'b0; 
    assign out[5320] = 1'b0; 
    assign out[5321] = 1'b0; 
    assign out[5322] = 1'b0; 
    assign out[5323] = 1'b0; 
    assign out[5324] = 1'b0; 
    assign out[5325] = 1'b0; 
    assign out[5326] = 1'b0; 
    assign out[5327] = 1'b0; 
    assign out[5328] = 1'b0; 
    assign out[5329] = 1'b0; 
    assign out[5330] = 1'b0; 
    assign out[5331] = 1'b0; 
    assign out[5332] = 1'b0; 
    assign out[5333] = 1'b0; 
    assign out[5334] = 1'b0; 
    assign out[5335] = 1'b0; 
    assign out[5336] = 1'b0; 
    assign out[5337] = 1'b0; 
    assign out[5338] = 1'b0; 
    assign out[5339] = 1'b0; 
    assign out[5340] = 1'b0; 
    assign out[5341] = 1'b0; 
    assign out[5342] = 1'b0; 
    assign out[5343] = 1'b0; 
    assign out[5344] = 1'b0; 
    assign out[5345] = 1'b0; 
    assign out[5346] = 1'b0; 
    assign out[5347] = 1'b0; 
    assign out[5348] = 1'b0; 
    assign out[5349] = 1'b0; 
    assign out[5350] = 1'b0; 
    assign out[5351] = 1'b0; 
    assign out[5352] = 1'b0; 
    assign out[5353] = 1'b0; 
    assign out[5354] = 1'b0; 
    assign out[5355] = 1'b0; 
    assign out[5356] = 1'b0; 
    assign out[5357] = 1'b0; 
    assign out[5358] = 1'b0; 
    assign out[5359] = 1'b0; 
    assign out[5360] = 1'b0; 
    assign out[5361] = 1'b0; 
    assign out[5362] = 1'b0; 
    assign out[5363] = 1'b0; 
    assign out[5364] = 1'b0; 
    assign out[5365] = 1'b0; 
    assign out[5366] = 1'b0; 
    assign out[5367] = 1'b0; 
    assign out[5368] = 1'b0; 
    assign out[5369] = 1'b0; 
    assign out[5370] = 1'b0; 
    assign out[5371] = 1'b0; 
    assign out[5372] = 1'b0; 
    assign out[5373] = 1'b0; 
    assign out[5374] = 1'b0; 
    assign out[5375] = 1'b0; 
    assign out[5376] = 1'b0; 
    assign out[5377] = 1'b0; 
    assign out[5378] = 1'b0; 
    assign out[5379] = 1'b0; 
    assign out[5380] = 1'b0; 
    assign out[5381] = 1'b0; 
    assign out[5382] = 1'b0; 
    assign out[5383] = 1'b0; 
    assign out[5384] = 1'b0; 
    assign out[5385] = 1'b0; 
    assign out[5386] = 1'b0; 
    assign out[5387] = 1'b0; 
    assign out[5388] = 1'b0; 
    assign out[5389] = 1'b0; 
    assign out[5390] = 1'b0; 
    assign out[5391] = 1'b0; 
    assign out[5392] = 1'b0; 
    assign out[5393] = 1'b0; 
    assign out[5394] = 1'b0; 
    assign out[5395] = 1'b0; 
    assign out[5396] = 1'b0; 
    assign out[5397] = 1'b0; 
    assign out[5398] = 1'b0; 
    assign out[5399] = 1'b0; 
    assign out[5400] = 1'b0; 
    assign out[5401] = 1'b0; 
    assign out[5402] = 1'b0; 
    assign out[5403] = 1'b0; 
    assign out[5404] = 1'b0; 
    assign out[5405] = 1'b0; 
    assign out[5406] = 1'b0; 
    assign out[5407] = 1'b0; 
    assign out[5408] = 1'b0; 
    assign out[5409] = 1'b0; 
    assign out[5410] = 1'b0; 
    assign out[5411] = 1'b0; 
    assign out[5412] = 1'b0; 
    assign out[5413] = 1'b0; 
    assign out[5414] = 1'b0; 
    assign out[5415] = 1'b0; 
    assign out[5416] = 1'b0; 
    assign out[5417] = 1'b0; 
    assign out[5418] = 1'b0; 
    assign out[5419] = 1'b0; 
    assign out[5420] = 1'b0; 
    assign out[5421] = 1'b0; 
    assign out[5422] = 1'b0; 
    assign out[5423] = 1'b0; 
    assign out[5424] = 1'b0; 
    assign out[5425] = 1'b0; 
    assign out[5426] = 1'b0; 
    assign out[5427] = 1'b0; 
    assign out[5428] = 1'b0; 
    assign out[5429] = 1'b0; 
    assign out[5430] = 1'b0; 
    assign out[5431] = 1'b0; 
    assign out[5432] = 1'b0; 
    assign out[5433] = 1'b0; 
    assign out[5434] = 1'b0; 
    assign out[5435] = 1'b0; 
    assign out[5436] = 1'b0; 
    assign out[5437] = 1'b0; 
    assign out[5438] = 1'b0; 
    assign out[5439] = 1'b0; 
    assign out[5440] = 1'b0; 
    assign out[5441] = 1'b0; 
    assign out[5442] = 1'b0; 
    assign out[5443] = 1'b0; 
    assign out[5444] = 1'b0; 
    assign out[5445] = 1'b0; 
    assign out[5446] = 1'b0; 
    assign out[5447] = 1'b0; 
    assign out[5448] = 1'b0; 
    assign out[5449] = 1'b0; 
    assign out[5450] = 1'b0; 
    assign out[5451] = 1'b0; 
    assign out[5452] = 1'b0; 
    assign out[5453] = 1'b0; 
    assign out[5454] = 1'b0; 
    assign out[5455] = 1'b0; 
    assign out[5456] = 1'b0; 
    assign out[5457] = 1'b0; 
    assign out[5458] = 1'b0; 
    assign out[5459] = 1'b0; 
    assign out[5460] = 1'b0; 
    assign out[5461] = 1'b0; 
    assign out[5462] = 1'b0; 
    assign out[5463] = 1'b0; 
    assign out[5464] = 1'b0; 
    assign out[5465] = 1'b0; 
    assign out[5466] = 1'b0; 
    assign out[5467] = 1'b0; 
    assign out[5468] = 1'b0; 
    assign out[5469] = 1'b0; 
    assign out[5470] = 1'b0; 
    assign out[5471] = 1'b0; 
    assign out[5472] = 1'b0; 
    assign out[5473] = 1'b0; 
    assign out[5474] = 1'b0; 
    assign out[5475] = 1'b0; 
    assign out[5476] = 1'b0; 
    assign out[5477] = 1'b0; 
    assign out[5478] = 1'b0; 
    assign out[5479] = 1'b0; 
    assign out[5480] = 1'b0; 
    assign out[5481] = 1'b0; 
    assign out[5482] = 1'b0; 
    assign out[5483] = 1'b0; 
    assign out[5484] = 1'b0; 
    assign out[5485] = 1'b0; 
    assign out[5486] = 1'b0; 
    assign out[5487] = 1'b0; 
    assign out[5488] = 1'b0; 
    assign out[5489] = 1'b0; 
    assign out[5490] = 1'b0; 
    assign out[5491] = 1'b0; 
    assign out[5492] = 1'b0; 
    assign out[5493] = 1'b0; 
    assign out[5494] = 1'b0; 
    assign out[5495] = 1'b0; 
    assign out[5496] = 1'b0; 
    assign out[5497] = 1'b0; 
    assign out[5498] = 1'b0; 
    assign out[5499] = 1'b0; 
    assign out[5500] = 1'b0; 
    assign out[5501] = 1'b0; 
    assign out[5502] = 1'b0; 
    assign out[5503] = 1'b0; 
    assign out[5504] = 1'b0; 
    assign out[5505] = 1'b0; 
    assign out[5506] = 1'b0; 
    assign out[5507] = 1'b0; 
    assign out[5508] = 1'b0; 
    assign out[5509] = 1'b0; 
    assign out[5510] = 1'b0; 
    assign out[5511] = 1'b0; 
    assign out[5512] = 1'b0; 
    assign out[5513] = 1'b0; 
    assign out[5514] = 1'b0; 
    assign out[5515] = 1'b0; 
    assign out[5516] = 1'b0; 
    assign out[5517] = 1'b0; 
    assign out[5518] = 1'b0; 
    assign out[5519] = 1'b0; 
    assign out[5520] = 1'b0; 
    assign out[5521] = 1'b0; 
    assign out[5522] = 1'b0; 
    assign out[5523] = 1'b0; 
    assign out[5524] = 1'b0; 
    assign out[5525] = 1'b0; 
    assign out[5526] = 1'b0; 
    assign out[5527] = 1'b0; 
    assign out[5528] = 1'b0; 
    assign out[5529] = 1'b0; 
    assign out[5530] = 1'b0; 
    assign out[5531] = 1'b0; 
    assign out[5532] = 1'b0; 
    assign out[5533] = 1'b0; 
    assign out[5534] = 1'b0; 
    assign out[5535] = 1'b0; 
    assign out[5536] = 1'b0; 
    assign out[5537] = 1'b0; 
    assign out[5538] = 1'b0; 
    assign out[5539] = 1'b0; 
    assign out[5540] = 1'b0; 
    assign out[5541] = 1'b0; 
    assign out[5542] = 1'b0; 
    assign out[5543] = 1'b0; 
    assign out[5544] = 1'b0; 
    assign out[5545] = 1'b0; 
    assign out[5546] = 1'b0; 
    assign out[5547] = 1'b0; 
    assign out[5548] = 1'b0; 
    assign out[5549] = 1'b0; 
    assign out[5550] = 1'b0; 
    assign out[5551] = 1'b0; 
    assign out[5552] = 1'b0; 
    assign out[5553] = 1'b0; 
    assign out[5554] = 1'b0; 
    assign out[5555] = 1'b0; 
    assign out[5556] = 1'b0; 
    assign out[5557] = 1'b0; 
    assign out[5558] = 1'b0; 
    assign out[5559] = 1'b0; 
    assign out[5560] = 1'b0; 
    assign out[5561] = 1'b0; 
    assign out[5562] = 1'b0; 
    assign out[5563] = 1'b0; 
    assign out[5564] = 1'b0; 
    assign out[5565] = 1'b0; 
    assign out[5566] = 1'b0; 
    assign out[5567] = 1'b0; 
    assign out[5568] = 1'b0; 
    assign out[5569] = 1'b0; 
    assign out[5570] = 1'b0; 
    assign out[5571] = 1'b0; 
    assign out[5572] = 1'b0; 
    assign out[5573] = 1'b0; 
    assign out[5574] = 1'b0; 
    assign out[5575] = 1'b0; 
    assign out[5576] = 1'b0; 
    assign out[5577] = 1'b0; 
    assign out[5578] = 1'b0; 
    assign out[5579] = 1'b0; 
    assign out[5580] = 1'b0; 
    assign out[5581] = 1'b0; 
    assign out[5582] = 1'b0; 
    assign out[5583] = 1'b0; 
    assign out[5584] = 1'b0; 
    assign out[5585] = 1'b0; 
    assign out[5586] = 1'b0; 
    assign out[5587] = 1'b0; 
    assign out[5588] = 1'b0; 
    assign out[5589] = 1'b0; 
    assign out[5590] = 1'b0; 
    assign out[5591] = 1'b0; 
    assign out[5592] = 1'b0; 
    assign out[5593] = 1'b0; 
    assign out[5594] = 1'b0; 
    assign out[5595] = 1'b0; 
    assign out[5596] = 1'b0; 
    assign out[5597] = 1'b0; 
    assign out[5598] = 1'b0; 
    assign out[5599] = 1'b0; 
    assign out[5600] = 1'b0; 
    assign out[5601] = 1'b0; 
    assign out[5602] = 1'b0; 
    assign out[5603] = 1'b0; 
    assign out[5604] = 1'b0; 
    assign out[5605] = 1'b0; 
    assign out[5606] = 1'b0; 
    assign out[5607] = 1'b0; 
    assign out[5608] = 1'b0; 
    assign out[5609] = 1'b0; 
    assign out[5610] = 1'b0; 
    assign out[5611] = 1'b0; 
    assign out[5612] = 1'b0; 
    assign out[5613] = 1'b0; 
    assign out[5614] = 1'b0; 
    assign out[5615] = 1'b0; 
    assign out[5616] = 1'b0; 
    assign out[5617] = 1'b0; 
    assign out[5618] = 1'b0; 
    assign out[5619] = 1'b0; 
    assign out[5620] = 1'b0; 
    assign out[5621] = 1'b0; 
    assign out[5622] = 1'b0; 
    assign out[5623] = 1'b0; 
    assign out[5624] = 1'b0; 
    assign out[5625] = 1'b0; 
    assign out[5626] = 1'b0; 
    assign out[5627] = 1'b0; 
    assign out[5628] = 1'b0; 
    assign out[5629] = 1'b0; 
    assign out[5630] = 1'b0; 
    assign out[5631] = 1'b0; 
    assign out[5632] = 1'b0; 
    assign out[5633] = 1'b0; 
    assign out[5634] = 1'b0; 
    assign out[5635] = 1'b0; 
    assign out[5636] = 1'b0; 
    assign out[5637] = 1'b0; 
    assign out[5638] = 1'b0; 
    assign out[5639] = 1'b0; 
    assign out[5640] = 1'b0; 
    assign out[5641] = 1'b0; 
    assign out[5642] = 1'b0; 
    assign out[5643] = 1'b0; 
    assign out[5644] = 1'b0; 
    assign out[5645] = 1'b0; 
    assign out[5646] = 1'b0; 
    assign out[5647] = 1'b0; 
    assign out[5648] = 1'b0; 
    assign out[5649] = 1'b0; 
    assign out[5650] = 1'b0; 
    assign out[5651] = 1'b0; 
    assign out[5652] = 1'b0; 
    assign out[5653] = 1'b0; 
    assign out[5654] = 1'b0; 
    assign out[5655] = 1'b0; 
    assign out[5656] = 1'b0; 
    assign out[5657] = 1'b0; 
    assign out[5658] = 1'b0; 
    assign out[5659] = 1'b0; 
    assign out[5660] = 1'b0; 
    assign out[5661] = 1'b0; 
    assign out[5662] = 1'b0; 
    assign out[5663] = 1'b0; 
    assign out[5664] = 1'b0; 
    assign out[5665] = 1'b0; 
    assign out[5666] = 1'b0; 
    assign out[5667] = 1'b0; 
    assign out[5668] = 1'b0; 
    assign out[5669] = 1'b0; 
    assign out[5670] = 1'b0; 
    assign out[5671] = 1'b0; 
    assign out[5672] = 1'b0; 
    assign out[5673] = 1'b0; 
    assign out[5674] = 1'b0; 
    assign out[5675] = 1'b0; 
    assign out[5676] = 1'b0; 
    assign out[5677] = 1'b0; 
    assign out[5678] = 1'b0; 
    assign out[5679] = 1'b0; 
    assign out[5680] = 1'b0; 
    assign out[5681] = 1'b0; 
    assign out[5682] = 1'b0; 
    assign out[5683] = 1'b0; 
    assign out[5684] = 1'b0; 
    assign out[5685] = 1'b0; 
    assign out[5686] = 1'b0; 
    assign out[5687] = 1'b0; 
    assign out[5688] = 1'b0; 
    assign out[5689] = 1'b0; 
    assign out[5690] = 1'b0; 
    assign out[5691] = 1'b0; 
    assign out[5692] = 1'b0; 
    assign out[5693] = 1'b0; 
    assign out[5694] = 1'b0; 
    assign out[5695] = 1'b0; 
    assign out[5696] = 1'b0; 
    assign out[5697] = 1'b0; 
    assign out[5698] = 1'b0; 
    assign out[5699] = 1'b0; 
    assign out[5700] = 1'b0; 
    assign out[5701] = 1'b0; 
    assign out[5702] = 1'b0; 
    assign out[5703] = 1'b0; 
    assign out[5704] = 1'b0; 
    assign out[5705] = 1'b0; 
    assign out[5706] = 1'b0; 
    assign out[5707] = 1'b0; 
    assign out[5708] = 1'b0; 
    assign out[5709] = 1'b0; 
    assign out[5710] = 1'b0; 
    assign out[5711] = 1'b0; 
    assign out[5712] = 1'b0; 
    assign out[5713] = 1'b0; 
    assign out[5714] = 1'b0; 
    assign out[5715] = 1'b0; 
    assign out[5716] = 1'b0; 
    assign out[5717] = 1'b0; 
    assign out[5718] = 1'b0; 
    assign out[5719] = 1'b0; 
    assign out[5720] = 1'b0; 
    assign out[5721] = 1'b0; 
    assign out[5722] = 1'b0; 
    assign out[5723] = 1'b0; 
    assign out[5724] = 1'b0; 
    assign out[5725] = 1'b0; 
    assign out[5726] = 1'b0; 
    assign out[5727] = 1'b0; 
    assign out[5728] = 1'b0; 
    assign out[5729] = 1'b0; 
    assign out[5730] = 1'b0; 
    assign out[5731] = 1'b0; 
    assign out[5732] = 1'b0; 
    assign out[5733] = 1'b0; 
    assign out[5734] = 1'b0; 
    assign out[5735] = 1'b0; 
    assign out[5736] = 1'b0; 
    assign out[5737] = 1'b0; 
    assign out[5738] = 1'b0; 
    assign out[5739] = 1'b0; 
    assign out[5740] = 1'b0; 
    assign out[5741] = 1'b0; 
    assign out[5742] = 1'b0; 
    assign out[5743] = 1'b0; 
    assign out[5744] = 1'b0; 
    assign out[5745] = 1'b0; 
    assign out[5746] = 1'b0; 
    assign out[5747] = 1'b0; 
    assign out[5748] = 1'b0; 
    assign out[5749] = 1'b0; 
    assign out[5750] = 1'b0; 
    assign out[5751] = 1'b0; 
    assign out[5752] = 1'b0; 
    assign out[5753] = 1'b0; 
    assign out[5754] = 1'b0; 
    assign out[5755] = 1'b0; 
    assign out[5756] = 1'b0; 
    assign out[5757] = 1'b0; 
    assign out[5758] = 1'b0; 
    assign out[5759] = 1'b0; 
    assign out[5760] = 1'b0; 
    assign out[5761] = 1'b0; 
    assign out[5762] = 1'b0; 
    assign out[5763] = 1'b0; 
    assign out[5764] = 1'b0; 
    assign out[5765] = 1'b0; 
    assign out[5766] = 1'b0; 
    assign out[5767] = 1'b0; 
    assign out[5768] = 1'b0; 
    assign out[5769] = 1'b0; 
    assign out[5770] = 1'b0; 
    assign out[5771] = 1'b0; 
    assign out[5772] = 1'b0; 
    assign out[5773] = 1'b0; 
    assign out[5774] = 1'b0; 
    assign out[5775] = 1'b0; 
    assign out[5776] = 1'b0; 
    assign out[5777] = 1'b0; 
    assign out[5778] = 1'b0; 
    assign out[5779] = 1'b0; 
    assign out[5780] = 1'b0; 
    assign out[5781] = 1'b0; 
    assign out[5782] = 1'b0; 
    assign out[5783] = 1'b0; 
    assign out[5784] = 1'b0; 
    assign out[5785] = 1'b0; 
    assign out[5786] = 1'b0; 
    assign out[5787] = 1'b0; 
    assign out[5788] = 1'b0; 
    assign out[5789] = 1'b0; 
    assign out[5790] = 1'b0; 
    assign out[5791] = 1'b0; 
    assign out[5792] = 1'b0; 
    assign out[5793] = 1'b0; 
    assign out[5794] = 1'b0; 
    assign out[5795] = 1'b0; 
    assign out[5796] = 1'b0; 
    assign out[5797] = 1'b0; 
    assign out[5798] = 1'b0; 
    assign out[5799] = 1'b0; 
    assign out[5800] = 1'b0; 
    assign out[5801] = 1'b0; 
    assign out[5802] = 1'b0; 
    assign out[5803] = 1'b0; 
    assign out[5804] = 1'b0; 
    assign out[5805] = 1'b0; 
    assign out[5806] = 1'b0; 
    assign out[5807] = 1'b0; 
    assign out[5808] = 1'b0; 
    assign out[5809] = 1'b0; 
    assign out[5810] = 1'b0; 
    assign out[5811] = 1'b0; 
    assign out[5812] = 1'b0; 
    assign out[5813] = 1'b0; 
    assign out[5814] = 1'b0; 
    assign out[5815] = 1'b0; 
    assign out[5816] = 1'b0; 
    assign out[5817] = 1'b0; 
    assign out[5818] = 1'b0; 
    assign out[5819] = 1'b0; 
    assign out[5820] = 1'b0; 
    assign out[5821] = 1'b0; 
    assign out[5822] = 1'b0; 
    assign out[5823] = 1'b0; 
    assign out[5824] = 1'b0; 
    assign out[5825] = 1'b0; 
    assign out[5826] = 1'b0; 
    assign out[5827] = 1'b0; 
    assign out[5828] = 1'b0; 
    assign out[5829] = 1'b0; 
    assign out[5830] = 1'b0; 
    assign out[5831] = 1'b0; 
    assign out[5832] = 1'b0; 
    assign out[5833] = 1'b0; 
    assign out[5834] = 1'b0; 
    assign out[5835] = 1'b0; 
    assign out[5836] = 1'b0; 
    assign out[5837] = 1'b0; 
    assign out[5838] = 1'b0; 
    assign out[5839] = 1'b0; 
    assign out[5840] = 1'b0; 
    assign out[5841] = 1'b0; 
    assign out[5842] = 1'b0; 
    assign out[5843] = 1'b0; 
    assign out[5844] = 1'b0; 
    assign out[5845] = 1'b0; 
    assign out[5846] = 1'b0; 
    assign out[5847] = 1'b0; 
    assign out[5848] = 1'b0; 
    assign out[5849] = 1'b0; 
    assign out[5850] = 1'b0; 
    assign out[5851] = 1'b0; 
    assign out[5852] = 1'b0; 
    assign out[5853] = 1'b0; 
    assign out[5854] = 1'b0; 
    assign out[5855] = 1'b0; 
    assign out[5856] = 1'b0; 
    assign out[5857] = 1'b0; 
    assign out[5858] = 1'b0; 
    assign out[5859] = 1'b0; 
    assign out[5860] = 1'b0; 
    assign out[5861] = 1'b0; 
    assign out[5862] = 1'b0; 
    assign out[5863] = 1'b0; 
    assign out[5864] = 1'b0; 
    assign out[5865] = 1'b0; 
    assign out[5866] = 1'b0; 
    assign out[5867] = 1'b0; 
    assign out[5868] = 1'b0; 
    assign out[5869] = 1'b0; 
    assign out[5870] = 1'b0; 
    assign out[5871] = 1'b0; 
    assign out[5872] = 1'b0; 
    assign out[5873] = 1'b0; 
    assign out[5874] = 1'b0; 
    assign out[5875] = 1'b0; 
    assign out[5876] = 1'b0; 
    assign out[5877] = 1'b0; 
    assign out[5878] = 1'b0; 
    assign out[5879] = 1'b0; 
    assign out[5880] = 1'b0; 
    assign out[5881] = 1'b0; 
    assign out[5882] = 1'b0; 
    assign out[5883] = 1'b0; 
    assign out[5884] = 1'b0; 
    assign out[5885] = 1'b0; 
    assign out[5886] = 1'b0; 
    assign out[5887] = 1'b0; 
    assign out[5888] = 1'b0; 
    assign out[5889] = 1'b0; 
    assign out[5890] = 1'b0; 
    assign out[5891] = 1'b0; 
    assign out[5892] = 1'b0; 
    assign out[5893] = 1'b0; 
    assign out[5894] = 1'b0; 
    assign out[5895] = 1'b0; 
    assign out[5896] = 1'b0; 
    assign out[5897] = 1'b0; 
    assign out[5898] = 1'b0; 
    assign out[5899] = 1'b0; 
    assign out[5900] = 1'b0; 
    assign out[5901] = 1'b0; 
    assign out[5902] = 1'b0; 
    assign out[5903] = 1'b0; 
    assign out[5904] = 1'b0; 
    assign out[5905] = 1'b0; 
    assign out[5906] = 1'b0; 
    assign out[5907] = 1'b0; 
    assign out[5908] = 1'b0; 
    assign out[5909] = 1'b0; 
    assign out[5910] = 1'b0; 
    assign out[5911] = 1'b0; 
    assign out[5912] = 1'b0; 
    assign out[5913] = 1'b0; 
    assign out[5914] = 1'b0; 
    assign out[5915] = 1'b0; 
    assign out[5916] = 1'b0; 
    assign out[5917] = 1'b0; 
    assign out[5918] = 1'b0; 
    assign out[5919] = 1'b0; 
    assign out[5920] = 1'b0; 
    assign out[5921] = 1'b0; 
    assign out[5922] = 1'b0; 
    assign out[5923] = 1'b0; 
    assign out[5924] = 1'b0; 
    assign out[5925] = 1'b0; 
    assign out[5926] = 1'b0; 
    assign out[5927] = 1'b0; 
    assign out[5928] = 1'b0; 
    assign out[5929] = 1'b0; 
    assign out[5930] = 1'b0; 
    assign out[5931] = 1'b0; 
    assign out[5932] = 1'b0; 
    assign out[5933] = 1'b0; 
    assign out[5934] = 1'b0; 
    assign out[5935] = 1'b0; 
    assign out[5936] = 1'b0; 
    assign out[5937] = 1'b0; 
    assign out[5938] = 1'b0; 
    assign out[5939] = 1'b0; 
    assign out[5940] = 1'b0; 
    assign out[5941] = 1'b0; 
    assign out[5942] = 1'b0; 
    assign out[5943] = 1'b0; 
    assign out[5944] = 1'b0; 
    assign out[5945] = 1'b0; 
    assign out[5946] = 1'b0; 
    assign out[5947] = 1'b0; 
    assign out[5948] = 1'b0; 
    assign out[5949] = 1'b0; 
    assign out[5950] = 1'b0; 
    assign out[5951] = 1'b0; 
    assign out[5952] = 1'b0; 
    assign out[5953] = 1'b0; 
    assign out[5954] = 1'b0; 
    assign out[5955] = 1'b0; 
    assign out[5956] = 1'b0; 
    assign out[5957] = 1'b0; 
    assign out[5958] = 1'b0; 
    assign out[5959] = 1'b0; 
    assign out[5960] = 1'b0; 
    assign out[5961] = 1'b0; 
    assign out[5962] = 1'b0; 
    assign out[5963] = 1'b0; 
    assign out[5964] = 1'b0; 
    assign out[5965] = 1'b0; 
    assign out[5966] = 1'b0; 
    assign out[5967] = 1'b0; 
    assign out[5968] = 1'b0; 
    assign out[5969] = 1'b0; 
    assign out[5970] = 1'b0; 
    assign out[5971] = 1'b0; 
    assign out[5972] = 1'b0; 
    assign out[5973] = 1'b0; 
    assign out[5974] = 1'b0; 
    assign out[5975] = 1'b0; 
    assign out[5976] = 1'b0; 
    assign out[5977] = 1'b0; 
    assign out[5978] = 1'b0; 
    assign out[5979] = 1'b0; 
    assign out[5980] = 1'b0; 
    assign out[5981] = 1'b0; 
    assign out[5982] = 1'b0; 
    assign out[5983] = 1'b0; 
    assign out[5984] = 1'b0; 
    assign out[5985] = 1'b0; 
    assign out[5986] = 1'b0; 
    assign out[5987] = 1'b0; 
    assign out[5988] = 1'b0; 
    assign out[5989] = 1'b0; 
    assign out[5990] = 1'b0; 
    assign out[5991] = 1'b0; 
    assign out[5992] = 1'b0; 
    assign out[5993] = 1'b0; 
    assign out[5994] = 1'b0; 
    assign out[5995] = 1'b0; 
    assign out[5996] = 1'b0; 
    assign out[5997] = 1'b0; 
    assign out[5998] = 1'b0; 
    assign out[5999] = 1'b0; 
    assign out[6000] = 1'b0; 
    assign out[6001] = 1'b0; 
    assign out[6002] = 1'b0; 
    assign out[6003] = 1'b0; 
    assign out[6004] = 1'b0; 
    assign out[6005] = 1'b0; 
    assign out[6006] = 1'b0; 
    assign out[6007] = 1'b0; 
    assign out[6008] = 1'b0; 
    assign out[6009] = 1'b0; 
    assign out[6010] = 1'b0; 
    assign out[6011] = 1'b0; 
    assign out[6012] = 1'b0; 
    assign out[6013] = 1'b0; 
    assign out[6014] = 1'b0; 
    assign out[6015] = 1'b0; 
    assign out[6016] = 1'b0; 
    assign out[6017] = 1'b0; 
    assign out[6018] = 1'b0; 
    assign out[6019] = 1'b0; 
    assign out[6020] = 1'b0; 
    assign out[6021] = 1'b0; 
    assign out[6022] = 1'b0; 
    assign out[6023] = 1'b0; 
    assign out[6024] = 1'b0; 
    assign out[6025] = 1'b0; 
    assign out[6026] = 1'b0; 
    assign out[6027] = 1'b0; 
    assign out[6028] = 1'b0; 
    assign out[6029] = 1'b0; 
    assign out[6030] = 1'b0; 
    assign out[6031] = 1'b0; 
    assign out[6032] = 1'b0; 
    assign out[6033] = 1'b0; 
    assign out[6034] = 1'b0; 
    assign out[6035] = 1'b0; 
    assign out[6036] = 1'b0; 
    assign out[6037] = 1'b0; 
    assign out[6038] = 1'b0; 
    assign out[6039] = 1'b0; 
    assign out[6040] = 1'b0; 
    assign out[6041] = 1'b0; 
    assign out[6042] = 1'b0; 
    assign out[6043] = 1'b0; 
    assign out[6044] = 1'b0; 
    assign out[6045] = 1'b0; 
    assign out[6046] = 1'b0; 
    assign out[6047] = 1'b0; 
    assign out[6048] = 1'b0; 
    assign out[6049] = 1'b0; 
    assign out[6050] = 1'b0; 
    assign out[6051] = 1'b0; 
    assign out[6052] = 1'b0; 
    assign out[6053] = 1'b0; 
    assign out[6054] = 1'b0; 
    assign out[6055] = 1'b0; 
    assign out[6056] = 1'b0; 
    assign out[6057] = 1'b0; 
    assign out[6058] = 1'b0; 
    assign out[6059] = 1'b0; 
    assign out[6060] = 1'b0; 
    assign out[6061] = 1'b0; 
    assign out[6062] = 1'b0; 
    assign out[6063] = 1'b0; 
    assign out[6064] = 1'b0; 
    assign out[6065] = 1'b0; 
    assign out[6066] = 1'b0; 
    assign out[6067] = 1'b0; 
    assign out[6068] = 1'b0; 
    assign out[6069] = 1'b0; 
    assign out[6070] = 1'b0; 
    assign out[6071] = 1'b0; 
    assign out[6072] = 1'b0; 
    assign out[6073] = 1'b0; 
    assign out[6074] = 1'b0; 
    assign out[6075] = 1'b0; 
    assign out[6076] = 1'b0; 
    assign out[6077] = 1'b0; 
    assign out[6078] = 1'b0; 
    assign out[6079] = 1'b0; 
    assign out[6080] = 1'b0; 
    assign out[6081] = 1'b0; 
    assign out[6082] = 1'b0; 
    assign out[6083] = 1'b0; 
    assign out[6084] = 1'b0; 
    assign out[6085] = 1'b0; 
    assign out[6086] = 1'b0; 
    assign out[6087] = 1'b0; 
    assign out[6088] = 1'b0; 
    assign out[6089] = 1'b0; 
    assign out[6090] = 1'b0; 
    assign out[6091] = 1'b0; 
    assign out[6092] = 1'b0; 
    assign out[6093] = 1'b0; 
    assign out[6094] = 1'b0; 
    assign out[6095] = 1'b0; 
    assign out[6096] = 1'b0; 
    assign out[6097] = 1'b0; 
    assign out[6098] = 1'b0; 
    assign out[6099] = 1'b0; 
    assign out[6100] = 1'b0; 
    assign out[6101] = 1'b0; 
    assign out[6102] = 1'b0; 
    assign out[6103] = 1'b0; 
    assign out[6104] = 1'b0; 
    assign out[6105] = 1'b0; 
    assign out[6106] = 1'b0; 
    assign out[6107] = 1'b0; 
    assign out[6108] = 1'b0; 
    assign out[6109] = 1'b0; 
    assign out[6110] = 1'b0; 
    assign out[6111] = 1'b0; 
    assign out[6112] = 1'b0; 
    assign out[6113] = 1'b0; 
    assign out[6114] = 1'b0; 
    assign out[6115] = 1'b0; 
    assign out[6116] = 1'b0; 
    assign out[6117] = 1'b0; 
    assign out[6118] = 1'b0; 
    assign out[6119] = 1'b0; 
    assign out[6120] = 1'b0; 
    assign out[6121] = 1'b0; 
    assign out[6122] = 1'b0; 
    assign out[6123] = 1'b0; 
    assign out[6124] = 1'b0; 
    assign out[6125] = 1'b0; 
    assign out[6126] = 1'b0; 
    assign out[6127] = 1'b0; 
    assign out[6128] = 1'b0; 
    assign out[6129] = 1'b0; 
    assign out[6130] = 1'b0; 
    assign out[6131] = 1'b0; 
    assign out[6132] = 1'b0; 
    assign out[6133] = 1'b0; 
    assign out[6134] = 1'b0; 
    assign out[6135] = 1'b0; 
    assign out[6136] = 1'b0; 
    assign out[6137] = 1'b0; 
    assign out[6138] = 1'b0; 
    assign out[6139] = 1'b0; 
    assign out[6140] = 1'b0; 
    assign out[6141] = 1'b0; 
    assign out[6142] = 1'b0; 
    assign out[6143] = 1'b0; 
    assign out[6144] = 1'b0; 
    assign out[6145] = 1'b0; 
    assign out[6146] = 1'b0; 
    assign out[6147] = 1'b0; 
    assign out[6148] = 1'b0; 
    assign out[6149] = 1'b0; 
    assign out[6150] = 1'b0; 
    assign out[6151] = 1'b0; 
    assign out[6152] = 1'b0; 
    assign out[6153] = 1'b0; 
    assign out[6154] = 1'b0; 
    assign out[6155] = 1'b0; 
    assign out[6156] = 1'b0; 
    assign out[6157] = 1'b0; 
    assign out[6158] = 1'b0; 
    assign out[6159] = 1'b0; 
    assign out[6160] = 1'b0; 
    assign out[6161] = 1'b0; 
    assign out[6162] = 1'b0; 
    assign out[6163] = 1'b0; 
    assign out[6164] = 1'b0; 
    assign out[6165] = 1'b0; 
    assign out[6166] = 1'b0; 
    assign out[6167] = 1'b0; 
    assign out[6168] = 1'b0; 
    assign out[6169] = 1'b0; 
    assign out[6170] = 1'b0; 
    assign out[6171] = 1'b0; 
    assign out[6172] = 1'b0; 
    assign out[6173] = 1'b0; 
    assign out[6174] = 1'b0; 
    assign out[6175] = 1'b0; 
    assign out[6176] = 1'b0; 
    assign out[6177] = 1'b0; 
    assign out[6178] = 1'b0; 
    assign out[6179] = 1'b0; 
    assign out[6180] = 1'b0; 
    assign out[6181] = 1'b0; 
    assign out[6182] = 1'b0; 
    assign out[6183] = 1'b0; 
    assign out[6184] = 1'b0; 
    assign out[6185] = 1'b0; 
    assign out[6186] = 1'b0; 
    assign out[6187] = 1'b0; 
    assign out[6188] = 1'b0; 
    assign out[6189] = 1'b0; 
    assign out[6190] = 1'b0; 
    assign out[6191] = 1'b0; 
    assign out[6192] = 1'b0; 
    assign out[6193] = 1'b0; 
    assign out[6194] = 1'b0; 
    assign out[6195] = 1'b0; 
    assign out[6196] = 1'b0; 
    assign out[6197] = 1'b0; 
    assign out[6198] = 1'b0; 
    assign out[6199] = 1'b0; 
    assign out[6200] = 1'b0; 
    assign out[6201] = 1'b0; 
    assign out[6202] = 1'b0; 
    assign out[6203] = 1'b0; 
    assign out[6204] = 1'b0; 
    assign out[6205] = 1'b0; 
    assign out[6206] = 1'b0; 
    assign out[6207] = 1'b0; 
    assign out[6208] = 1'b0; 
    assign out[6209] = 1'b0; 
    assign out[6210] = 1'b0; 
    assign out[6211] = 1'b0; 
    assign out[6212] = 1'b0; 
    assign out[6213] = 1'b0; 
    assign out[6214] = 1'b0; 
    assign out[6215] = 1'b0; 
    assign out[6216] = 1'b0; 
    assign out[6217] = 1'b0; 
    assign out[6218] = 1'b0; 
    assign out[6219] = 1'b0; 
    assign out[6220] = 1'b0; 
    assign out[6221] = 1'b0; 
    assign out[6222] = 1'b0; 
    assign out[6223] = 1'b0; 
    assign out[6224] = 1'b0; 
    assign out[6225] = 1'b0; 
    assign out[6226] = 1'b0; 
    assign out[6227] = 1'b0; 
    assign out[6228] = 1'b0; 
    assign out[6229] = 1'b0; 
    assign out[6230] = 1'b0; 
    assign out[6231] = 1'b0; 
    assign out[6232] = 1'b0; 
    assign out[6233] = 1'b0; 
    assign out[6234] = 1'b0; 
    assign out[6235] = 1'b0; 
    assign out[6236] = 1'b0; 
    assign out[6237] = 1'b0; 
    assign out[6238] = 1'b0; 
    assign out[6239] = 1'b0; 
    assign out[6240] = 1'b0; 
    assign out[6241] = 1'b0; 
    assign out[6242] = 1'b0; 
    assign out[6243] = 1'b0; 
    assign out[6244] = 1'b0; 
    assign out[6245] = 1'b0; 
    assign out[6246] = 1'b0; 
    assign out[6247] = 1'b0; 
    assign out[6248] = 1'b0; 
    assign out[6249] = 1'b0; 
    assign out[6250] = 1'b0; 
    assign out[6251] = 1'b0; 
    assign out[6252] = 1'b0; 
    assign out[6253] = 1'b0; 
    assign out[6254] = 1'b0; 
    assign out[6255] = 1'b0; 
    assign out[6256] = 1'b0; 
    assign out[6257] = 1'b0; 
    assign out[6258] = 1'b0; 
    assign out[6259] = 1'b0; 
    assign out[6260] = 1'b0; 
    assign out[6261] = 1'b0; 
    assign out[6262] = 1'b0; 
    assign out[6263] = 1'b0; 
    assign out[6264] = 1'b0; 
    assign out[6265] = 1'b0; 
    assign out[6266] = 1'b0; 
    assign out[6267] = 1'b0; 
    assign out[6268] = 1'b0; 
    assign out[6269] = 1'b0; 
    assign out[6270] = 1'b0; 
    assign out[6271] = 1'b0; 
    assign out[6272] = 1'b0; 
    assign out[6273] = 1'b0; 
    assign out[6274] = 1'b0; 
    assign out[6275] = 1'b0; 
    assign out[6276] = 1'b0; 
    assign out[6277] = 1'b0; 
    assign out[6278] = 1'b0; 
    assign out[6279] = 1'b0; 
    assign out[6280] = 1'b0; 
    assign out[6281] = 1'b0; 
    assign out[6282] = 1'b0; 
    assign out[6283] = 1'b0; 
    assign out[6284] = 1'b0; 
    assign out[6285] = 1'b0; 
    assign out[6286] = 1'b0; 
    assign out[6287] = 1'b0; 
    assign out[6288] = 1'b0; 
    assign out[6289] = 1'b0; 
    assign out[6290] = 1'b0; 
    assign out[6291] = 1'b0; 
    assign out[6292] = 1'b0; 
    assign out[6293] = 1'b0; 
    assign out[6294] = 1'b0; 
    assign out[6295] = 1'b0; 
    assign out[6296] = 1'b0; 
    assign out[6297] = 1'b0; 
    assign out[6298] = 1'b0; 
    assign out[6299] = 1'b0; 
    assign out[6300] = 1'b0; 
    assign out[6301] = 1'b0; 
    assign out[6302] = 1'b0; 
    assign out[6303] = 1'b0; 
    assign out[6304] = 1'b0; 
    assign out[6305] = 1'b0; 
    assign out[6306] = 1'b0; 
    assign out[6307] = 1'b0; 
    assign out[6308] = 1'b0; 
    assign out[6309] = 1'b0; 
    assign out[6310] = 1'b0; 
    assign out[6311] = 1'b0; 
    assign out[6312] = 1'b0; 
    assign out[6313] = 1'b0; 
    assign out[6314] = 1'b0; 
    assign out[6315] = 1'b0; 
    assign out[6316] = 1'b0; 
    assign out[6317] = 1'b0; 
    assign out[6318] = 1'b0; 
    assign out[6319] = 1'b0; 
    assign out[6320] = 1'b0; 
    assign out[6321] = 1'b0; 
    assign out[6322] = 1'b0; 
    assign out[6323] = 1'b0; 
    assign out[6324] = 1'b0; 
    assign out[6325] = 1'b0; 
    assign out[6326] = 1'b0; 
    assign out[6327] = 1'b0; 
    assign out[6328] = 1'b0; 
    assign out[6329] = 1'b0; 
    assign out[6330] = 1'b0; 
    assign out[6331] = 1'b0; 
    assign out[6332] = 1'b0; 
    assign out[6333] = 1'b0; 
    assign out[6334] = 1'b0; 
    assign out[6335] = 1'b0; 
    assign out[6336] = 1'b0; 
    assign out[6337] = 1'b0; 
    assign out[6338] = 1'b0; 
    assign out[6339] = 1'b0; 
    assign out[6340] = 1'b0; 
    assign out[6341] = 1'b0; 
    assign out[6342] = 1'b0; 
    assign out[6343] = 1'b0; 
    assign out[6344] = 1'b0; 
    assign out[6345] = 1'b0; 
    assign out[6346] = 1'b0; 
    assign out[6347] = 1'b0; 
    assign out[6348] = 1'b0; 
    assign out[6349] = 1'b0; 
    assign out[6350] = 1'b0; 
    assign out[6351] = 1'b0; 
    assign out[6352] = 1'b0; 
    assign out[6353] = 1'b0; 
    assign out[6354] = 1'b0; 
    assign out[6355] = 1'b0; 
    assign out[6356] = 1'b0; 
    assign out[6357] = 1'b0; 
    assign out[6358] = 1'b0; 
    assign out[6359] = 1'b0; 
    assign out[6360] = 1'b0; 
    assign out[6361] = 1'b0; 
    assign out[6362] = 1'b0; 
    assign out[6363] = 1'b0; 
    assign out[6364] = 1'b0; 
    assign out[6365] = 1'b0; 
    assign out[6366] = 1'b0; 
    assign out[6367] = 1'b0; 
    assign out[6368] = 1'b0; 
    assign out[6369] = 1'b0; 
    assign out[6370] = 1'b0; 
    assign out[6371] = 1'b0; 
    assign out[6372] = 1'b0; 
    assign out[6373] = 1'b0; 
    assign out[6374] = 1'b0; 
    assign out[6375] = 1'b0; 
    assign out[6376] = 1'b0; 
    assign out[6377] = 1'b0; 
    assign out[6378] = 1'b0; 
    assign out[6379] = 1'b0; 
    assign out[6380] = 1'b0; 
    assign out[6381] = 1'b0; 
    assign out[6382] = 1'b0; 
    assign out[6383] = 1'b0; 
    assign out[6384] = 1'b0; 
    assign out[6385] = 1'b0; 
    assign out[6386] = 1'b0; 
    assign out[6387] = 1'b0; 
    assign out[6388] = 1'b0; 
    assign out[6389] = 1'b0; 
    assign out[6390] = 1'b0; 
    assign out[6391] = 1'b0; 
    assign out[6392] = 1'b0; 
    assign out[6393] = 1'b0; 
    assign out[6394] = 1'b0; 
    assign out[6395] = 1'b0; 
    assign out[6396] = 1'b0; 
    assign out[6397] = 1'b0; 
    assign out[6398] = 1'b0; 
    assign out[6399] = 1'b0; 
    assign out[6400] = 1'b0; 
    assign out[6401] = 1'b0; 
    assign out[6402] = 1'b0; 
    assign out[6403] = 1'b0; 
    assign out[6404] = 1'b0; 
    assign out[6405] = 1'b0; 
    assign out[6406] = 1'b0; 
    assign out[6407] = 1'b0; 
    assign out[6408] = 1'b0; 
    assign out[6409] = 1'b0; 
    assign out[6410] = 1'b0; 
    assign out[6411] = 1'b0; 
    assign out[6412] = 1'b0; 
    assign out[6413] = 1'b0; 
    assign out[6414] = 1'b0; 
    assign out[6415] = 1'b0; 
    assign out[6416] = 1'b0; 
    assign out[6417] = 1'b0; 
    assign out[6418] = 1'b0; 
    assign out[6419] = 1'b0; 
    assign out[6420] = 1'b0; 
    assign out[6421] = 1'b0; 
    assign out[6422] = 1'b0; 
    assign out[6423] = 1'b0; 
    assign out[6424] = 1'b0; 
    assign out[6425] = 1'b0; 
    assign out[6426] = 1'b0; 
    assign out[6427] = 1'b0; 
    assign out[6428] = 1'b0; 
    assign out[6429] = 1'b0; 
    assign out[6430] = 1'b0; 
    assign out[6431] = 1'b0; 
    assign out[6432] = 1'b0; 
    assign out[6433] = 1'b0; 
    assign out[6434] = 1'b0; 
    assign out[6435] = 1'b0; 
    assign out[6436] = 1'b0; 
    assign out[6437] = 1'b0; 
    assign out[6438] = 1'b0; 
    assign out[6439] = 1'b0; 
    assign out[6440] = 1'b0; 
    assign out[6441] = 1'b0; 
    assign out[6442] = 1'b0; 
    assign out[6443] = 1'b0; 
    assign out[6444] = 1'b0; 
    assign out[6445] = 1'b0; 
    assign out[6446] = 1'b0; 
    assign out[6447] = 1'b0; 
    assign out[6448] = 1'b0; 
    assign out[6449] = 1'b0; 
    assign out[6450] = 1'b0; 
    assign out[6451] = 1'b0; 
    assign out[6452] = 1'b0; 
    assign out[6453] = 1'b0; 
    assign out[6454] = 1'b0; 
    assign out[6455] = 1'b0; 
    assign out[6456] = 1'b0; 
    assign out[6457] = 1'b0; 
    assign out[6458] = 1'b0; 
    assign out[6459] = 1'b0; 
    assign out[6460] = 1'b0; 
    assign out[6461] = 1'b0; 
    assign out[6462] = 1'b0; 
    assign out[6463] = 1'b0; 
    assign out[6464] = 1'b0; 
    assign out[6465] = 1'b0; 
    assign out[6466] = 1'b0; 
    assign out[6467] = 1'b0; 
    assign out[6468] = 1'b0; 
    assign out[6469] = 1'b0; 
    assign out[6470] = 1'b0; 
    assign out[6471] = 1'b0; 
    assign out[6472] = 1'b0; 
    assign out[6473] = 1'b0; 
    assign out[6474] = 1'b0; 
    assign out[6475] = 1'b0; 
    assign out[6476] = 1'b0; 
    assign out[6477] = 1'b0; 
    assign out[6478] = 1'b0; 
    assign out[6479] = 1'b0; 
    assign out[6480] = 1'b0; 
    assign out[6481] = 1'b0; 
    assign out[6482] = 1'b0; 
    assign out[6483] = 1'b0; 
    assign out[6484] = 1'b0; 
    assign out[6485] = 1'b0; 
    assign out[6486] = 1'b0; 
    assign out[6487] = 1'b0; 
    assign out[6488] = 1'b0; 
    assign out[6489] = 1'b0; 
    assign out[6490] = 1'b0; 
    assign out[6491] = 1'b0; 
    assign out[6492] = 1'b0; 
    assign out[6493] = 1'b0; 
    assign out[6494] = 1'b0; 
    assign out[6495] = 1'b0; 
    assign out[6496] = 1'b0; 
    assign out[6497] = 1'b0; 
    assign out[6498] = 1'b0; 
    assign out[6499] = 1'b0; 
    assign out[6500] = 1'b0; 
    assign out[6501] = 1'b0; 
    assign out[6502] = 1'b0; 
    assign out[6503] = 1'b0; 
    assign out[6504] = 1'b0; 
    assign out[6505] = 1'b0; 
    assign out[6506] = 1'b0; 
    assign out[6507] = 1'b0; 
    assign out[6508] = 1'b0; 
    assign out[6509] = 1'b0; 
    assign out[6510] = 1'b0; 
    assign out[6511] = 1'b0; 
    assign out[6512] = 1'b0; 
    assign out[6513] = 1'b0; 
    assign out[6514] = 1'b0; 
    assign out[6515] = 1'b0; 
    assign out[6516] = 1'b0; 
    assign out[6517] = 1'b0; 
    assign out[6518] = 1'b0; 
    assign out[6519] = 1'b0; 
    assign out[6520] = 1'b0; 
    assign out[6521] = 1'b0; 
    assign out[6522] = 1'b0; 
    assign out[6523] = 1'b0; 
    assign out[6524] = 1'b0; 
    assign out[6525] = 1'b0; 
    assign out[6526] = 1'b0; 
    assign out[6527] = 1'b0; 
    assign out[6528] = 1'b0; 
    assign out[6529] = 1'b0; 
    assign out[6530] = 1'b0; 
    assign out[6531] = 1'b0; 
    assign out[6532] = 1'b0; 
    assign out[6533] = 1'b0; 
    assign out[6534] = 1'b0; 
    assign out[6535] = 1'b0; 
    assign out[6536] = 1'b0; 
    assign out[6537] = 1'b0; 
    assign out[6538] = 1'b0; 
    assign out[6539] = 1'b0; 
    assign out[6540] = 1'b0; 
    assign out[6541] = 1'b0; 
    assign out[6542] = 1'b0; 
    assign out[6543] = 1'b0; 
    assign out[6544] = 1'b0; 
    assign out[6545] = 1'b0; 
    assign out[6546] = 1'b0; 
    assign out[6547] = 1'b0; 
    assign out[6548] = 1'b0; 
    assign out[6549] = 1'b0; 
    assign out[6550] = 1'b0; 
    assign out[6551] = 1'b0; 
    assign out[6552] = 1'b0; 
    assign out[6553] = 1'b0; 
    assign out[6554] = 1'b0; 
    assign out[6555] = 1'b0; 
    assign out[6556] = 1'b0; 
    assign out[6557] = 1'b0; 
    assign out[6558] = 1'b0; 
    assign out[6559] = 1'b0; 
    assign out[6560] = 1'b0; 
    assign out[6561] = 1'b0; 
    assign out[6562] = 1'b0; 
    assign out[6563] = 1'b0; 
    assign out[6564] = 1'b0; 
    assign out[6565] = 1'b0; 
    assign out[6566] = 1'b0; 
    assign out[6567] = 1'b0; 
    assign out[6568] = 1'b0; 
    assign out[6569] = 1'b0; 
    assign out[6570] = 1'b0; 
    assign out[6571] = 1'b0; 
    assign out[6572] = 1'b0; 
    assign out[6573] = 1'b0; 
    assign out[6574] = 1'b0; 
    assign out[6575] = 1'b0; 
    assign out[6576] = 1'b0; 
    assign out[6577] = 1'b0; 
    assign out[6578] = 1'b0; 
    assign out[6579] = 1'b0; 
    assign out[6580] = 1'b0; 
    assign out[6581] = 1'b0; 
    assign out[6582] = 1'b0; 
    assign out[6583] = 1'b0; 
    assign out[6584] = 1'b0; 
    assign out[6585] = 1'b0; 
    assign out[6586] = 1'b0; 
    assign out[6587] = 1'b0; 
    assign out[6588] = 1'b0; 
    assign out[6589] = 1'b0; 
    assign out[6590] = 1'b0; 
    assign out[6591] = 1'b0; 
    assign out[6592] = 1'b0; 
    assign out[6593] = 1'b0; 
    assign out[6594] = 1'b0; 
    assign out[6595] = 1'b0; 
    assign out[6596] = 1'b0; 
    assign out[6597] = 1'b0; 
    assign out[6598] = 1'b0; 
    assign out[6599] = 1'b0; 
    assign out[6600] = 1'b0; 
    assign out[6601] = 1'b0; 
    assign out[6602] = 1'b0; 
    assign out[6603] = 1'b0; 
    assign out[6604] = 1'b0; 
    assign out[6605] = 1'b0; 
    assign out[6606] = 1'b0; 
    assign out[6607] = 1'b0; 
    assign out[6608] = 1'b0; 
    assign out[6609] = 1'b0; 
    assign out[6610] = 1'b0; 
    assign out[6611] = 1'b0; 
    assign out[6612] = 1'b0; 
    assign out[6613] = 1'b0; 
    assign out[6614] = 1'b0; 
    assign out[6615] = 1'b0; 
    assign out[6616] = 1'b0; 
    assign out[6617] = 1'b0; 
    assign out[6618] = 1'b0; 
    assign out[6619] = 1'b0; 
    assign out[6620] = 1'b0; 
    assign out[6621] = 1'b0; 
    assign out[6622] = 1'b0; 
    assign out[6623] = 1'b0; 
    assign out[6624] = 1'b0; 
    assign out[6625] = 1'b0; 
    assign out[6626] = 1'b0; 
    assign out[6627] = 1'b0; 
    assign out[6628] = 1'b0; 
    assign out[6629] = 1'b0; 
    assign out[6630] = 1'b0; 
    assign out[6631] = 1'b0; 
    assign out[6632] = 1'b0; 
    assign out[6633] = 1'b0; 
    assign out[6634] = 1'b0; 
    assign out[6635] = 1'b0; 
    assign out[6636] = 1'b0; 
    assign out[6637] = 1'b0; 
    assign out[6638] = 1'b0; 
    assign out[6639] = 1'b0; 
    assign out[6640] = 1'b0; 
    assign out[6641] = 1'b0; 
    assign out[6642] = 1'b0; 
    assign out[6643] = 1'b0; 
    assign out[6644] = 1'b0; 
    assign out[6645] = 1'b0; 
    assign out[6646] = 1'b0; 
    assign out[6647] = 1'b0; 
    assign out[6648] = 1'b0; 
    assign out[6649] = 1'b0; 
    assign out[6650] = 1'b0; 
    assign out[6651] = 1'b0; 
    assign out[6652] = 1'b0; 
    assign out[6653] = 1'b0; 
    assign out[6654] = 1'b0; 
    assign out[6655] = 1'b0; 
    assign out[6656] = 1'b0; 
    assign out[6657] = 1'b0; 
    assign out[6658] = 1'b0; 
    assign out[6659] = 1'b0; 
    assign out[6660] = 1'b0; 
    assign out[6661] = 1'b0; 
    assign out[6662] = 1'b0; 
    assign out[6663] = 1'b0; 
    assign out[6664] = 1'b0; 
    assign out[6665] = 1'b0; 
    assign out[6666] = 1'b0; 
    assign out[6667] = 1'b0; 
    assign out[6668] = 1'b0; 
    assign out[6669] = 1'b0; 
    assign out[6670] = 1'b0; 
    assign out[6671] = 1'b0; 
    assign out[6672] = 1'b0; 
    assign out[6673] = 1'b0; 
    assign out[6674] = 1'b0; 
    assign out[6675] = 1'b0; 
    assign out[6676] = 1'b0; 
    assign out[6677] = 1'b0; 
    assign out[6678] = 1'b0; 
    assign out[6679] = 1'b0; 
    assign out[6680] = 1'b0; 
    assign out[6681] = 1'b0; 
    assign out[6682] = 1'b0; 
    assign out[6683] = 1'b0; 
    assign out[6684] = 1'b0; 
    assign out[6685] = 1'b0; 
    assign out[6686] = 1'b0; 
    assign out[6687] = 1'b0; 
    assign out[6688] = 1'b0; 
    assign out[6689] = 1'b0; 
    assign out[6690] = 1'b0; 
    assign out[6691] = 1'b0; 
    assign out[6692] = 1'b0; 
    assign out[6693] = 1'b0; 
    assign out[6694] = 1'b0; 
    assign out[6695] = 1'b0; 
    assign out[6696] = 1'b0; 
    assign out[6697] = 1'b0; 
    assign out[6698] = 1'b0; 
    assign out[6699] = 1'b0; 
    assign out[6700] = 1'b0; 
    assign out[6701] = 1'b0; 
    assign out[6702] = 1'b0; 
    assign out[6703] = 1'b0; 
    assign out[6704] = 1'b0; 
    assign out[6705] = 1'b0; 
    assign out[6706] = 1'b0; 
    assign out[6707] = 1'b0; 
    assign out[6708] = 1'b0; 
    assign out[6709] = 1'b0; 
    assign out[6710] = 1'b0; 
    assign out[6711] = 1'b0; 
    assign out[6712] = 1'b0; 
    assign out[6713] = 1'b0; 
    assign out[6714] = 1'b0; 
    assign out[6715] = 1'b0; 
    assign out[6716] = 1'b0; 
    assign out[6717] = 1'b0; 
    assign out[6718] = 1'b0; 
    assign out[6719] = 1'b0; 
    assign out[6720] = 1'b0; 
    assign out[6721] = 1'b0; 
    assign out[6722] = 1'b0; 
    assign out[6723] = 1'b0; 
    assign out[6724] = 1'b0; 
    assign out[6725] = 1'b0; 
    assign out[6726] = 1'b0; 
    assign out[6727] = 1'b0; 
    assign out[6728] = 1'b0; 
    assign out[6729] = 1'b0; 
    assign out[6730] = 1'b0; 
    assign out[6731] = 1'b0; 
    assign out[6732] = 1'b0; 
    assign out[6733] = 1'b0; 
    assign out[6734] = 1'b0; 
    assign out[6735] = 1'b0; 
    assign out[6736] = 1'b0; 
    assign out[6737] = 1'b0; 
    assign out[6738] = 1'b0; 
    assign out[6739] = 1'b0; 
    assign out[6740] = 1'b0; 
    assign out[6741] = 1'b0; 
    assign out[6742] = 1'b0; 
    assign out[6743] = 1'b0; 
    assign out[6744] = 1'b0; 
    assign out[6745] = 1'b0; 
    assign out[6746] = 1'b0; 
    assign out[6747] = 1'b0; 
    assign out[6748] = 1'b0; 
    assign out[6749] = 1'b0; 
    assign out[6750] = 1'b0; 
    assign out[6751] = 1'b0; 
    assign out[6752] = 1'b0; 
    assign out[6753] = 1'b0; 
    assign out[6754] = 1'b0; 
    assign out[6755] = 1'b0; 
    assign out[6756] = 1'b0; 
    assign out[6757] = 1'b0; 
    assign out[6758] = 1'b0; 
    assign out[6759] = 1'b0; 
    assign out[6760] = 1'b0; 
    assign out[6761] = 1'b0; 
    assign out[6762] = 1'b0; 
    assign out[6763] = 1'b0; 
    assign out[6764] = 1'b0; 
    assign out[6765] = 1'b0; 
    assign out[6766] = 1'b0; 
    assign out[6767] = 1'b0; 
    assign out[6768] = 1'b0; 
    assign out[6769] = 1'b0; 
    assign out[6770] = 1'b0; 
    assign out[6771] = 1'b0; 
    assign out[6772] = 1'b0; 
    assign out[6773] = 1'b0; 
    assign out[6774] = 1'b0; 
    assign out[6775] = 1'b0; 
    assign out[6776] = 1'b0; 
    assign out[6777] = 1'b0; 
    assign out[6778] = 1'b0; 
    assign out[6779] = 1'b0; 
    assign out[6780] = 1'b0; 
    assign out[6781] = 1'b0; 
    assign out[6782] = 1'b0; 
    assign out[6783] = 1'b0; 
    assign out[6784] = 1'b0; 
    assign out[6785] = 1'b0; 
    assign out[6786] = 1'b0; 
    assign out[6787] = 1'b0; 
    assign out[6788] = 1'b0; 
    assign out[6789] = 1'b0; 
    assign out[6790] = 1'b0; 
    assign out[6791] = 1'b0; 
    assign out[6792] = 1'b0; 
    assign out[6793] = 1'b0; 
    assign out[6794] = 1'b0; 
    assign out[6795] = 1'b0; 
    assign out[6796] = 1'b0; 
    assign out[6797] = 1'b0; 
    assign out[6798] = 1'b0; 
    assign out[6799] = 1'b0; 
    assign out[6800] = 1'b0; 
    assign out[6801] = 1'b0; 
    assign out[6802] = 1'b0; 
    assign out[6803] = 1'b0; 
    assign out[6804] = 1'b0; 
    assign out[6805] = 1'b0; 
    assign out[6806] = 1'b0; 
    assign out[6807] = 1'b0; 
    assign out[6808] = 1'b0; 
    assign out[6809] = 1'b0; 
    assign out[6810] = 1'b0; 
    assign out[6811] = 1'b0; 
    assign out[6812] = 1'b0; 
    assign out[6813] = 1'b0; 
    assign out[6814] = 1'b0; 
    assign out[6815] = 1'b0; 
    assign out[6816] = 1'b0; 
    assign out[6817] = 1'b0; 
    assign out[6818] = 1'b0; 
    assign out[6819] = 1'b0; 
    assign out[6820] = 1'b0; 
    assign out[6821] = 1'b0; 
    assign out[6822] = 1'b0; 
    assign out[6823] = 1'b0; 
    assign out[6824] = 1'b0; 
    assign out[6825] = 1'b0; 
    assign out[6826] = 1'b0; 
    assign out[6827] = 1'b0; 
    assign out[6828] = 1'b0; 
    assign out[6829] = 1'b0; 
    assign out[6830] = 1'b0; 
    assign out[6831] = 1'b0; 
    assign out[6832] = 1'b0; 
    assign out[6833] = 1'b0; 
    assign out[6834] = 1'b0; 
    assign out[6835] = 1'b0; 
    assign out[6836] = 1'b0; 
    assign out[6837] = 1'b0; 
    assign out[6838] = 1'b0; 
    assign out[6839] = 1'b0; 
    assign out[6840] = 1'b0; 
    assign out[6841] = 1'b0; 
    assign out[6842] = 1'b0; 
    assign out[6843] = 1'b0; 
    assign out[6844] = 1'b0; 
    assign out[6845] = 1'b0; 
    assign out[6846] = 1'b0; 
    assign out[6847] = 1'b0; 
    assign out[6848] = 1'b0; 
    assign out[6849] = 1'b0; 
    assign out[6850] = 1'b0; 
    assign out[6851] = 1'b0; 
    assign out[6852] = 1'b0; 
    assign out[6853] = 1'b0; 
    assign out[6854] = 1'b0; 
    assign out[6855] = 1'b0; 
    assign out[6856] = 1'b0; 
    assign out[6857] = 1'b0; 
    assign out[6858] = 1'b0; 
    assign out[6859] = 1'b0; 
    assign out[6860] = 1'b0; 
    assign out[6861] = 1'b0; 
    assign out[6862] = 1'b0; 
    assign out[6863] = 1'b0; 
    assign out[6864] = 1'b0; 
    assign out[6865] = 1'b0; 
    assign out[6866] = 1'b0; 
    assign out[6867] = 1'b0; 
    assign out[6868] = 1'b0; 
    assign out[6869] = 1'b0; 
    assign out[6870] = 1'b0; 
    assign out[6871] = 1'b0; 
    assign out[6872] = 1'b0; 
    assign out[6873] = 1'b0; 
    assign out[6874] = 1'b0; 
    assign out[6875] = 1'b0; 
    assign out[6876] = 1'b0; 
    assign out[6877] = 1'b0; 
    assign out[6878] = 1'b0; 
    assign out[6879] = 1'b0; 
    assign out[6880] = 1'b0; 
    assign out[6881] = 1'b0; 
    assign out[6882] = 1'b0; 
    assign out[6883] = 1'b0; 
    assign out[6884] = 1'b0; 
    assign out[6885] = 1'b0; 
    assign out[6886] = 1'b0; 
    assign out[6887] = 1'b0; 
    assign out[6888] = 1'b0; 
    assign out[6889] = 1'b0; 
    assign out[6890] = 1'b0; 
    assign out[6891] = 1'b0; 
    assign out[6892] = 1'b0; 
    assign out[6893] = 1'b0; 
    assign out[6894] = 1'b0; 
    assign out[6895] = 1'b0; 
    assign out[6896] = 1'b0; 
    assign out[6897] = 1'b0; 
    assign out[6898] = 1'b0; 
    assign out[6899] = 1'b0; 
    assign out[6900] = 1'b0; 
    assign out[6901] = 1'b0; 
    assign out[6902] = 1'b0; 
    assign out[6903] = 1'b0; 
    assign out[6904] = 1'b0; 
    assign out[6905] = 1'b0; 
    assign out[6906] = 1'b0; 
    assign out[6907] = 1'b0; 
    assign out[6908] = 1'b0; 
    assign out[6909] = 1'b0; 
    assign out[6910] = 1'b0; 
    assign out[6911] = 1'b0; 
    assign out[6912] = 1'b0; 
    assign out[6913] = 1'b0; 
    assign out[6914] = 1'b0; 
    assign out[6915] = 1'b0; 
    assign out[6916] = 1'b0; 
    assign out[6917] = 1'b0; 
    assign out[6918] = 1'b0; 
    assign out[6919] = 1'b0; 
    assign out[6920] = 1'b0; 
    assign out[6921] = 1'b0; 
    assign out[6922] = 1'b0; 
    assign out[6923] = 1'b0; 
    assign out[6924] = 1'b0; 
    assign out[6925] = 1'b0; 
    assign out[6926] = 1'b0; 
    assign out[6927] = 1'b0; 
    assign out[6928] = 1'b0; 
    assign out[6929] = 1'b0; 
    assign out[6930] = 1'b0; 
    assign out[6931] = 1'b0; 
    assign out[6932] = 1'b0; 
    assign out[6933] = 1'b0; 
    assign out[6934] = 1'b0; 
    assign out[6935] = 1'b0; 
    assign out[6936] = 1'b0; 
    assign out[6937] = 1'b0; 
    assign out[6938] = 1'b0; 
    assign out[6939] = 1'b0; 
    assign out[6940] = 1'b0; 
    assign out[6941] = 1'b0; 
    assign out[6942] = 1'b0; 
    assign out[6943] = 1'b0; 
    assign out[6944] = 1'b0; 
    assign out[6945] = 1'b0; 
    assign out[6946] = 1'b0; 
    assign out[6947] = 1'b0; 
    assign out[6948] = 1'b0; 
    assign out[6949] = 1'b0; 
    assign out[6950] = 1'b0; 
    assign out[6951] = 1'b0; 
    assign out[6952] = 1'b0; 
    assign out[6953] = 1'b0; 
    assign out[6954] = 1'b0; 
    assign out[6955] = 1'b0; 
    assign out[6956] = 1'b0; 
    assign out[6957] = 1'b0; 
    assign out[6958] = 1'b0; 
    assign out[6959] = 1'b0; 
    assign out[6960] = 1'b0; 
    assign out[6961] = 1'b0; 
    assign out[6962] = 1'b0; 
    assign out[6963] = 1'b0; 
    assign out[6964] = 1'b0; 
    assign out[6965] = 1'b0; 
    assign out[6966] = 1'b0; 
    assign out[6967] = 1'b0; 
    assign out[6968] = 1'b0; 
    assign out[6969] = 1'b0; 
    assign out[6970] = 1'b0; 
    assign out[6971] = 1'b0; 
    assign out[6972] = 1'b0; 
    assign out[6973] = 1'b0; 
    assign out[6974] = 1'b0; 
    assign out[6975] = 1'b0; 
    assign out[6976] = 1'b0; 
    assign out[6977] = 1'b0; 
    assign out[6978] = 1'b0; 
    assign out[6979] = 1'b0; 
    assign out[6980] = 1'b0; 
    assign out[6981] = 1'b0; 
    assign out[6982] = 1'b0; 
    assign out[6983] = 1'b0; 
    assign out[6984] = 1'b0; 
    assign out[6985] = 1'b0; 
    assign out[6986] = 1'b0; 
    assign out[6987] = 1'b0; 
    assign out[6988] = 1'b0; 
    assign out[6989] = 1'b0; 
    assign out[6990] = 1'b0; 
    assign out[6991] = 1'b0; 
    assign out[6992] = 1'b0; 
    assign out[6993] = 1'b0; 
    assign out[6994] = 1'b0; 
    assign out[6995] = 1'b0; 
    assign out[6996] = 1'b0; 
    assign out[6997] = 1'b0; 
    assign out[6998] = 1'b0; 
    assign out[6999] = 1'b0; 
    assign out[7000] = 1'b0; 
    assign out[7001] = 1'b0; 
    assign out[7002] = 1'b0; 
    assign out[7003] = 1'b0; 
    assign out[7004] = 1'b0; 
    assign out[7005] = 1'b0; 
    assign out[7006] = 1'b0; 
    assign out[7007] = 1'b0; 
    assign out[7008] = 1'b0; 
    assign out[7009] = 1'b0; 
    assign out[7010] = 1'b0; 
    assign out[7011] = 1'b0; 
    assign out[7012] = 1'b0; 
    assign out[7013] = 1'b0; 
    assign out[7014] = 1'b0; 
    assign out[7015] = 1'b0; 
    assign out[7016] = 1'b0; 
    assign out[7017] = 1'b0; 
    assign out[7018] = 1'b0; 
    assign out[7019] = 1'b0; 
    assign out[7020] = 1'b0; 
    assign out[7021] = 1'b0; 
    assign out[7022] = 1'b0; 
    assign out[7023] = 1'b0; 
    assign out[7024] = 1'b0; 
    assign out[7025] = 1'b0; 
    assign out[7026] = 1'b0; 
    assign out[7027] = 1'b0; 
    assign out[7028] = 1'b0; 
    assign out[7029] = 1'b0; 
    assign out[7030] = 1'b0; 
    assign out[7031] = 1'b0; 
    assign out[7032] = 1'b0; 
    assign out[7033] = 1'b0; 
    assign out[7034] = 1'b0; 
    assign out[7035] = 1'b0; 
    assign out[7036] = 1'b0; 
    assign out[7037] = 1'b0; 
    assign out[7038] = 1'b0; 
    assign out[7039] = 1'b0; 
    assign out[7040] = 1'b0; 
    assign out[7041] = 1'b0; 
    assign out[7042] = 1'b0; 
    assign out[7043] = 1'b0; 
    assign out[7044] = 1'b0; 
    assign out[7045] = 1'b0; 
    assign out[7046] = 1'b0; 
    assign out[7047] = 1'b0; 
    assign out[7048] = 1'b0; 
    assign out[7049] = 1'b0; 
    assign out[7050] = 1'b0; 
    assign out[7051] = 1'b0; 
    assign out[7052] = 1'b0; 
    assign out[7053] = 1'b0; 
    assign out[7054] = 1'b0; 
    assign out[7055] = 1'b0; 
    assign out[7056] = 1'b0; 
    assign out[7057] = 1'b0; 
    assign out[7058] = 1'b0; 
    assign out[7059] = 1'b0; 
    assign out[7060] = 1'b0; 
    assign out[7061] = 1'b0; 
    assign out[7062] = 1'b0; 
    assign out[7063] = 1'b0; 
    assign out[7064] = 1'b0; 
    assign out[7065] = 1'b0; 
    assign out[7066] = 1'b0; 
    assign out[7067] = 1'b0; 
    assign out[7068] = 1'b0; 
    assign out[7069] = 1'b0; 
    assign out[7070] = 1'b0; 
    assign out[7071] = 1'b0; 
    assign out[7072] = 1'b0; 
    assign out[7073] = 1'b0; 
    assign out[7074] = 1'b0; 
    assign out[7075] = 1'b0; 
    assign out[7076] = 1'b0; 
    assign out[7077] = 1'b0; 
    assign out[7078] = 1'b0; 
    assign out[7079] = 1'b0; 
    assign out[7080] = 1'b0; 
    assign out[7081] = 1'b0; 
    assign out[7082] = 1'b0; 
    assign out[7083] = 1'b0; 
    assign out[7084] = 1'b0; 
    assign out[7085] = 1'b0; 
    assign out[7086] = 1'b0; 
    assign out[7087] = 1'b0; 
    assign out[7088] = 1'b0; 
    assign out[7089] = 1'b0; 
    assign out[7090] = 1'b0; 
    assign out[7091] = 1'b0; 
    assign out[7092] = 1'b0; 
    assign out[7093] = 1'b0; 
    assign out[7094] = 1'b0; 
    assign out[7095] = 1'b0; 
    assign out[7096] = 1'b0; 
    assign out[7097] = 1'b0; 
    assign out[7098] = 1'b0; 
    assign out[7099] = 1'b0; 
    assign out[7100] = 1'b0; 
    assign out[7101] = 1'b0; 
    assign out[7102] = 1'b0; 
    assign out[7103] = 1'b0; 
    assign out[7104] = 1'b0; 
    assign out[7105] = 1'b0; 
    assign out[7106] = 1'b0; 
    assign out[7107] = 1'b0; 
    assign out[7108] = 1'b0; 
    assign out[7109] = 1'b0; 
    assign out[7110] = 1'b0; 
    assign out[7111] = 1'b0; 
    assign out[7112] = 1'b0; 
    assign out[7113] = 1'b0; 
    assign out[7114] = 1'b0; 
    assign out[7115] = 1'b0; 
    assign out[7116] = 1'b0; 
    assign out[7117] = 1'b0; 
    assign out[7118] = 1'b0; 
    assign out[7119] = 1'b0; 
    assign out[7120] = 1'b0; 
    assign out[7121] = 1'b0; 
    assign out[7122] = 1'b0; 
    assign out[7123] = 1'b0; 
    assign out[7124] = 1'b0; 
    assign out[7125] = 1'b0; 
    assign out[7126] = 1'b0; 
    assign out[7127] = 1'b0; 
    assign out[7128] = 1'b0; 
    assign out[7129] = 1'b0; 
    assign out[7130] = 1'b0; 
    assign out[7131] = 1'b0; 
    assign out[7132] = 1'b0; 
    assign out[7133] = 1'b0; 
    assign out[7134] = 1'b0; 
    assign out[7135] = 1'b0; 
    assign out[7136] = 1'b0; 
    assign out[7137] = 1'b0; 
    assign out[7138] = 1'b0; 
    assign out[7139] = 1'b0; 
    assign out[7140] = 1'b0; 
    assign out[7141] = 1'b0; 
    assign out[7142] = 1'b0; 
    assign out[7143] = 1'b0; 
    assign out[7144] = 1'b0; 
    assign out[7145] = 1'b0; 
    assign out[7146] = 1'b0; 
    assign out[7147] = 1'b0; 
    assign out[7148] = 1'b0; 
    assign out[7149] = 1'b0; 
    assign out[7150] = 1'b0; 
    assign out[7151] = 1'b0; 
    assign out[7152] = 1'b0; 
    assign out[7153] = 1'b0; 
    assign out[7154] = 1'b0; 
    assign out[7155] = 1'b0; 
    assign out[7156] = 1'b0; 
    assign out[7157] = 1'b0; 
    assign out[7158] = 1'b0; 
    assign out[7159] = 1'b0; 
    assign out[7160] = 1'b0; 
    assign out[7161] = 1'b0; 
    assign out[7162] = 1'b0; 
    assign out[7163] = 1'b0; 
    assign out[7164] = 1'b0; 
    assign out[7165] = 1'b0; 
    assign out[7166] = 1'b0; 
    assign out[7167] = 1'b0; 
    assign out[7168] = 1'b0; 
    assign out[7169] = 1'b0; 
    assign out[7170] = 1'b0; 
    assign out[7171] = 1'b0; 
    assign out[7172] = 1'b0; 
    assign out[7173] = 1'b0; 
    assign out[7174] = 1'b0; 
    assign out[7175] = 1'b0; 
    assign out[7176] = 1'b0; 
    assign out[7177] = 1'b0; 
    assign out[7178] = 1'b0; 
    assign out[7179] = 1'b0; 
    assign out[7180] = 1'b0; 
    assign out[7181] = 1'b0; 
    assign out[7182] = 1'b0; 
    assign out[7183] = 1'b0; 
    assign out[7184] = 1'b0; 
    assign out[7185] = 1'b0; 
    assign out[7186] = 1'b0; 
    assign out[7187] = 1'b0; 
    assign out[7188] = 1'b0; 
    assign out[7189] = 1'b0; 
    assign out[7190] = 1'b0; 
    assign out[7191] = 1'b0; 
    assign out[7192] = 1'b0; 
    assign out[7193] = 1'b0; 
    assign out[7194] = 1'b0; 
    assign out[7195] = 1'b0; 
    assign out[7196] = 1'b0; 
    assign out[7197] = 1'b0; 
    assign out[7198] = 1'b0; 
    assign out[7199] = 1'b0; 
    assign out[7200] = 1'b0; 
    assign out[7201] = 1'b0; 
    assign out[7202] = 1'b0; 
    assign out[7203] = 1'b0; 
    assign out[7204] = 1'b0; 
    assign out[7205] = 1'b0; 
    assign out[7206] = 1'b0; 
    assign out[7207] = 1'b0; 
    assign out[7208] = 1'b0; 
    assign out[7209] = 1'b0; 
    assign out[7210] = 1'b0; 
    assign out[7211] = 1'b0; 
    assign out[7212] = 1'b0; 
    assign out[7213] = 1'b0; 
    assign out[7214] = 1'b0; 
    assign out[7215] = 1'b0; 
    assign out[7216] = 1'b0; 
    assign out[7217] = 1'b0; 
    assign out[7218] = 1'b0; 
    assign out[7219] = 1'b0; 
    assign out[7220] = 1'b0; 
    assign out[7221] = 1'b0; 
    assign out[7222] = 1'b0; 
    assign out[7223] = 1'b0; 
    assign out[7224] = 1'b0; 
    assign out[7225] = 1'b0; 
    assign out[7226] = 1'b0; 
    assign out[7227] = 1'b0; 
    assign out[7228] = 1'b0; 
    assign out[7229] = 1'b0; 
    assign out[7230] = 1'b0; 
    assign out[7231] = 1'b0; 
    assign out[7232] = 1'b0; 
    assign out[7233] = 1'b0; 
    assign out[7234] = 1'b0; 
    assign out[7235] = 1'b0; 
    assign out[7236] = 1'b0; 
    assign out[7237] = 1'b0; 
    assign out[7238] = 1'b0; 
    assign out[7239] = 1'b0; 
    assign out[7240] = 1'b0; 
    assign out[7241] = 1'b0; 
    assign out[7242] = 1'b0; 
    assign out[7243] = 1'b0; 
    assign out[7244] = 1'b0; 
    assign out[7245] = 1'b0; 
    assign out[7246] = 1'b0; 
    assign out[7247] = 1'b0; 
    assign out[7248] = 1'b0; 
    assign out[7249] = 1'b0; 
    assign out[7250] = 1'b0; 
    assign out[7251] = 1'b0; 
    assign out[7252] = 1'b0; 
    assign out[7253] = 1'b0; 
    assign out[7254] = 1'b0; 
    assign out[7255] = 1'b0; 
    assign out[7256] = 1'b0; 
    assign out[7257] = 1'b0; 
    assign out[7258] = 1'b0; 
    assign out[7259] = 1'b0; 
    assign out[7260] = 1'b0; 
    assign out[7261] = 1'b0; 
    assign out[7262] = 1'b0; 
    assign out[7263] = 1'b0; 
    assign out[7264] = 1'b0; 
    assign out[7265] = 1'b0; 
    assign out[7266] = 1'b0; 
    assign out[7267] = 1'b0; 
    assign out[7268] = 1'b0; 
    assign out[7269] = 1'b0; 
    assign out[7270] = 1'b0; 
    assign out[7271] = 1'b0; 
    assign out[7272] = 1'b0; 
    assign out[7273] = 1'b0; 
    assign out[7274] = 1'b0; 
    assign out[7275] = 1'b0; 
    assign out[7276] = 1'b0; 
    assign out[7277] = 1'b0; 
    assign out[7278] = 1'b0; 
    assign out[7279] = 1'b0; 
    assign out[7280] = 1'b0; 
    assign out[7281] = 1'b0; 
    assign out[7282] = 1'b0; 
    assign out[7283] = 1'b0; 
    assign out[7284] = 1'b0; 
    assign out[7285] = 1'b0; 
    assign out[7286] = 1'b0; 
    assign out[7287] = 1'b0; 
    assign out[7288] = 1'b0; 
    assign out[7289] = 1'b0; 
    assign out[7290] = 1'b0; 
    assign out[7291] = 1'b0; 
    assign out[7292] = 1'b0; 
    assign out[7293] = 1'b0; 
    assign out[7294] = 1'b0; 
    assign out[7295] = 1'b0; 
    assign out[7296] = 1'b0; 
    assign out[7297] = 1'b0; 
    assign out[7298] = 1'b0; 
    assign out[7299] = 1'b0; 
    assign out[7300] = 1'b0; 
    assign out[7301] = 1'b0; 
    assign out[7302] = 1'b0; 
    assign out[7303] = 1'b0; 
    assign out[7304] = 1'b0; 
    assign out[7305] = 1'b0; 
    assign out[7306] = 1'b0; 
    assign out[7307] = 1'b0; 
    assign out[7308] = 1'b0; 
    assign out[7309] = 1'b0; 
    assign out[7310] = 1'b0; 
    assign out[7311] = 1'b0; 
    assign out[7312] = 1'b0; 
    assign out[7313] = 1'b0; 
    assign out[7314] = 1'b0; 
    assign out[7315] = 1'b0; 
    assign out[7316] = 1'b0; 
    assign out[7317] = 1'b0; 
    assign out[7318] = 1'b0; 
    assign out[7319] = 1'b0; 
    assign out[7320] = 1'b0; 
    assign out[7321] = 1'b0; 
    assign out[7322] = 1'b0; 
    assign out[7323] = 1'b0; 
    assign out[7324] = 1'b0; 
    assign out[7325] = 1'b0; 
    assign out[7326] = 1'b0; 
    assign out[7327] = 1'b0; 
    assign out[7328] = 1'b0; 
    assign out[7329] = 1'b0; 
    assign out[7330] = 1'b0; 
    assign out[7331] = 1'b0; 
    assign out[7332] = 1'b0; 
    assign out[7333] = 1'b0; 
    assign out[7334] = 1'b0; 
    assign out[7335] = 1'b0; 
    assign out[7336] = 1'b0; 
    assign out[7337] = 1'b0; 
    assign out[7338] = 1'b0; 
    assign out[7339] = 1'b0; 
    assign out[7340] = 1'b0; 
    assign out[7341] = 1'b0; 
    assign out[7342] = 1'b0; 
    assign out[7343] = 1'b0; 
    assign out[7344] = 1'b0; 
    assign out[7345] = 1'b0; 
    assign out[7346] = 1'b0; 
    assign out[7347] = 1'b0; 
    assign out[7348] = 1'b0; 
    assign out[7349] = 1'b0; 
    assign out[7350] = 1'b0; 
    assign out[7351] = 1'b0; 
    assign out[7352] = 1'b0; 
    assign out[7353] = 1'b0; 
    assign out[7354] = 1'b0; 
    assign out[7355] = 1'b0; 
    assign out[7356] = 1'b0; 
    assign out[7357] = 1'b0; 
    assign out[7358] = 1'b0; 
    assign out[7359] = 1'b0; 
    assign out[7360] = 1'b0; 
    assign out[7361] = 1'b0; 
    assign out[7362] = 1'b0; 
    assign out[7363] = 1'b0; 
    assign out[7364] = 1'b0; 
    assign out[7365] = 1'b0; 
    assign out[7366] = 1'b0; 
    assign out[7367] = 1'b0; 
    assign out[7368] = 1'b0; 
    assign out[7369] = 1'b0; 
    assign out[7370] = 1'b0; 
    assign out[7371] = 1'b0; 
    assign out[7372] = 1'b0; 
    assign out[7373] = 1'b0; 
    assign out[7374] = 1'b0; 
    assign out[7375] = 1'b0; 
    assign out[7376] = 1'b0; 
    assign out[7377] = 1'b0; 
    assign out[7378] = 1'b0; 
    assign out[7379] = 1'b0; 
    assign out[7380] = 1'b0; 
    assign out[7381] = 1'b0; 
    assign out[7382] = 1'b0; 
    assign out[7383] = 1'b0; 
    assign out[7384] = 1'b0; 
    assign out[7385] = 1'b0; 
    assign out[7386] = 1'b0; 
    assign out[7387] = 1'b0; 
    assign out[7388] = 1'b0; 
    assign out[7389] = 1'b0; 
    assign out[7390] = 1'b0; 
    assign out[7391] = 1'b0; 
    assign out[7392] = 1'b0; 
    assign out[7393] = 1'b0; 
    assign out[7394] = 1'b0; 
    assign out[7395] = 1'b0; 
    assign out[7396] = 1'b0; 
    assign out[7397] = 1'b0; 
    assign out[7398] = 1'b0; 
    assign out[7399] = 1'b0; 
    assign out[7400] = 1'b0; 
    assign out[7401] = 1'b0; 
    assign out[7402] = 1'b0; 
    assign out[7403] = 1'b0; 
    assign out[7404] = 1'b0; 
    assign out[7405] = 1'b0; 
    assign out[7406] = 1'b0; 
    assign out[7407] = 1'b0; 
    assign out[7408] = 1'b0; 
    assign out[7409] = 1'b0; 
    assign out[7410] = 1'b0; 
    assign out[7411] = 1'b0; 
    assign out[7412] = 1'b0; 
    assign out[7413] = 1'b0; 
    assign out[7414] = 1'b0; 
    assign out[7415] = 1'b0; 
    assign out[7416] = 1'b0; 
    assign out[7417] = 1'b0; 
    assign out[7418] = 1'b0; 
    assign out[7419] = 1'b0; 
    assign out[7420] = 1'b0; 
    assign out[7421] = 1'b0; 
    assign out[7422] = 1'b0; 
    assign out[7423] = 1'b0; 
    assign out[7424] = 1'b0; 
    assign out[7425] = 1'b0; 
    assign out[7426] = 1'b0; 
    assign out[7427] = 1'b0; 
    assign out[7428] = 1'b0; 
    assign out[7429] = 1'b0; 
    assign out[7430] = 1'b0; 
    assign out[7431] = 1'b0; 
    assign out[7432] = 1'b0; 
    assign out[7433] = 1'b0; 
    assign out[7434] = 1'b0; 
    assign out[7435] = 1'b0; 
    assign out[7436] = 1'b0; 
    assign out[7437] = 1'b0; 
    assign out[7438] = 1'b0; 
    assign out[7439] = 1'b0; 
    assign out[7440] = 1'b0; 
    assign out[7441] = 1'b0; 
    assign out[7442] = 1'b0; 
    assign out[7443] = 1'b0; 
    assign out[7444] = 1'b0; 
    assign out[7445] = 1'b0; 
    assign out[7446] = 1'b0; 
    assign out[7447] = 1'b0; 
    assign out[7448] = 1'b0; 
    assign out[7449] = 1'b0; 
    assign out[7450] = 1'b0; 
    assign out[7451] = 1'b0; 
    assign out[7452] = 1'b0; 
    assign out[7453] = 1'b0; 
    assign out[7454] = 1'b0; 
    assign out[7455] = 1'b0; 
    assign out[7456] = 1'b0; 
    assign out[7457] = 1'b0; 
    assign out[7458] = 1'b0; 
    assign out[7459] = 1'b0; 
    assign out[7460] = 1'b0; 
    assign out[7461] = 1'b0; 
    assign out[7462] = 1'b0; 
    assign out[7463] = 1'b0; 
    assign out[7464] = 1'b0; 
    assign out[7465] = 1'b0; 
    assign out[7466] = 1'b0; 
    assign out[7467] = 1'b0; 
    assign out[7468] = 1'b0; 
    assign out[7469] = 1'b0; 
    assign out[7470] = 1'b0; 
    assign out[7471] = 1'b0; 
    assign out[7472] = 1'b0; 
    assign out[7473] = 1'b0; 
    assign out[7474] = 1'b0; 
    assign out[7475] = 1'b0; 
    assign out[7476] = 1'b0; 
    assign out[7477] = 1'b0; 
    assign out[7478] = 1'b0; 
    assign out[7479] = 1'b0; 
    assign out[7480] = 1'b0; 
    assign out[7481] = 1'b0; 
    assign out[7482] = 1'b0; 
    assign out[7483] = 1'b0; 
    assign out[7484] = 1'b0; 
    assign out[7485] = 1'b0; 
    assign out[7486] = 1'b0; 
    assign out[7487] = 1'b0; 
    assign out[7488] = 1'b0; 
    assign out[7489] = 1'b0; 
    assign out[7490] = 1'b0; 
    assign out[7491] = 1'b0; 
    assign out[7492] = 1'b0; 
    assign out[7493] = 1'b0; 
    assign out[7494] = 1'b0; 
    assign out[7495] = 1'b0; 
    assign out[7496] = 1'b0; 
    assign out[7497] = 1'b0; 
    assign out[7498] = 1'b0; 
    assign out[7499] = 1'b0; 
    assign out[7500] = 1'b0; 
    assign out[7501] = 1'b0; 
    assign out[7502] = 1'b0; 
    assign out[7503] = 1'b0; 
    assign out[7504] = 1'b0; 
    assign out[7505] = 1'b0; 
    assign out[7506] = 1'b0; 
    assign out[7507] = 1'b0; 
    assign out[7508] = 1'b0; 
    assign out[7509] = 1'b0; 
    assign out[7510] = 1'b0; 
    assign out[7511] = 1'b0; 
    assign out[7512] = 1'b0; 
    assign out[7513] = 1'b0; 
    assign out[7514] = 1'b0; 
    assign out[7515] = 1'b0; 
    assign out[7516] = 1'b0; 
    assign out[7517] = 1'b0; 
    assign out[7518] = 1'b0; 
    assign out[7519] = 1'b0; 
    assign out[7520] = 1'b0; 
    assign out[7521] = 1'b0; 
    assign out[7522] = 1'b0; 
    assign out[7523] = 1'b0; 
    assign out[7524] = 1'b0; 
    assign out[7525] = 1'b0; 
    assign out[7526] = 1'b0; 
    assign out[7527] = 1'b0; 
    assign out[7528] = 1'b0; 
    assign out[7529] = 1'b0; 
    assign out[7530] = 1'b0; 
    assign out[7531] = 1'b0; 
    assign out[7532] = 1'b0; 
    assign out[7533] = 1'b0; 
    assign out[7534] = 1'b0; 
    assign out[7535] = 1'b0; 
    assign out[7536] = 1'b0; 
    assign out[7537] = 1'b0; 
    assign out[7538] = 1'b0; 
    assign out[7539] = 1'b0; 
    assign out[7540] = 1'b0; 
    assign out[7541] = 1'b0; 
    assign out[7542] = 1'b0; 
    assign out[7543] = 1'b0; 
    assign out[7544] = 1'b0; 
    assign out[7545] = 1'b0; 
    assign out[7546] = 1'b0; 
    assign out[7547] = 1'b0; 
    assign out[7548] = 1'b0; 
    assign out[7549] = 1'b0; 
    assign out[7550] = 1'b0; 
    assign out[7551] = 1'b0; 
    assign out[7552] = 1'b0; 
    assign out[7553] = 1'b0; 
    assign out[7554] = 1'b0; 
    assign out[7555] = 1'b0; 
    assign out[7556] = 1'b0; 
    assign out[7557] = 1'b0; 
    assign out[7558] = 1'b0; 
    assign out[7559] = 1'b0; 
    assign out[7560] = 1'b0; 
    assign out[7561] = 1'b0; 
    assign out[7562] = 1'b0; 
    assign out[7563] = 1'b0; 
    assign out[7564] = 1'b0; 
    assign out[7565] = 1'b0; 
    assign out[7566] = 1'b0; 
    assign out[7567] = 1'b0; 
    assign out[7568] = 1'b0; 
    assign out[7569] = 1'b0; 
    assign out[7570] = 1'b0; 
    assign out[7571] = 1'b0; 
    assign out[7572] = 1'b0; 
    assign out[7573] = 1'b0; 
    assign out[7574] = 1'b0; 
    assign out[7575] = 1'b0; 
    assign out[7576] = 1'b0; 
    assign out[7577] = 1'b0; 
    assign out[7578] = 1'b0; 
    assign out[7579] = 1'b0; 
    assign out[7580] = 1'b0; 
    assign out[7581] = 1'b0; 
    assign out[7582] = 1'b0; 
    assign out[7583] = 1'b0; 
    assign out[7584] = 1'b0; 
    assign out[7585] = 1'b0; 
    assign out[7586] = 1'b0; 
    assign out[7587] = 1'b0; 
    assign out[7588] = 1'b0; 
    assign out[7589] = 1'b0; 
    assign out[7590] = 1'b0; 
    assign out[7591] = 1'b0; 
    assign out[7592] = 1'b0; 
    assign out[7593] = 1'b0; 
    assign out[7594] = 1'b0; 
    assign out[7595] = 1'b0; 
    assign out[7596] = 1'b0; 
    assign out[7597] = 1'b0; 
    assign out[7598] = 1'b0; 
    assign out[7599] = 1'b0; 
    assign out[7600] = 1'b0; 
    assign out[7601] = 1'b0; 
    assign out[7602] = 1'b0; 
    assign out[7603] = 1'b0; 
    assign out[7604] = 1'b0; 
    assign out[7605] = 1'b0; 
    assign out[7606] = 1'b0; 
    assign out[7607] = 1'b0; 
    assign out[7608] = 1'b0; 
    assign out[7609] = 1'b0; 
    assign out[7610] = 1'b0; 
    assign out[7611] = 1'b0; 
    assign out[7612] = 1'b0; 
    assign out[7613] = 1'b0; 
    assign out[7614] = 1'b0; 
    assign out[7615] = 1'b0; 
    assign out[7616] = 1'b0; 
    assign out[7617] = 1'b0; 
    assign out[7618] = 1'b0; 
    assign out[7619] = 1'b0; 
    assign out[7620] = 1'b0; 
    assign out[7621] = 1'b0; 
    assign out[7622] = 1'b0; 
    assign out[7623] = 1'b0; 
    assign out[7624] = 1'b0; 
    assign out[7625] = 1'b0; 
    assign out[7626] = 1'b0; 
    assign out[7627] = 1'b0; 
    assign out[7628] = 1'b0; 
    assign out[7629] = 1'b0; 
    assign out[7630] = 1'b0; 
    assign out[7631] = 1'b0; 
    assign out[7632] = 1'b0; 
    assign out[7633] = 1'b0; 
    assign out[7634] = 1'b0; 
    assign out[7635] = 1'b0; 
    assign out[7636] = 1'b0; 
    assign out[7637] = 1'b0; 
    assign out[7638] = 1'b0; 
    assign out[7639] = 1'b0; 
    assign out[7640] = 1'b0; 
    assign out[7641] = 1'b0; 
    assign out[7642] = 1'b0; 
    assign out[7643] = 1'b0; 
    assign out[7644] = 1'b0; 
    assign out[7645] = 1'b0; 
    assign out[7646] = 1'b0; 
    assign out[7647] = 1'b0; 
    assign out[7648] = 1'b0; 
    assign out[7649] = 1'b0; 
    assign out[7650] = 1'b0; 
    assign out[7651] = 1'b0; 
    assign out[7652] = 1'b0; 
    assign out[7653] = 1'b0; 
    assign out[7654] = 1'b0; 
    assign out[7655] = 1'b0; 
    assign out[7656] = 1'b0; 
    assign out[7657] = 1'b0; 
    assign out[7658] = 1'b0; 
    assign out[7659] = 1'b0; 
    assign out[7660] = 1'b0; 
    assign out[7661] = 1'b0; 
    assign out[7662] = 1'b0; 
    assign out[7663] = 1'b0; 
    assign out[7664] = 1'b0; 
    assign out[7665] = 1'b0; 
    assign out[7666] = 1'b0; 
    assign out[7667] = 1'b0; 
    assign out[7668] = 1'b0; 
    assign out[7669] = 1'b0; 
    assign out[7670] = 1'b0; 
    assign out[7671] = 1'b0; 
    assign out[7672] = 1'b0; 
    assign out[7673] = 1'b0; 
    assign out[7674] = 1'b0; 
    assign out[7675] = 1'b0; 
    assign out[7676] = 1'b0; 
    assign out[7677] = 1'b0; 
    assign out[7678] = 1'b0; 
    assign out[7679] = 1'b0; 
    assign out[7680] = 1'b0; 
    assign out[7681] = 1'b0; 
    assign out[7682] = 1'b0; 
    assign out[7683] = 1'b0; 
    assign out[7684] = 1'b0; 
    assign out[7685] = 1'b0; 
    assign out[7686] = 1'b0; 
    assign out[7687] = 1'b0; 
    assign out[7688] = 1'b0; 
    assign out[7689] = 1'b0; 
    assign out[7690] = 1'b0; 
    assign out[7691] = 1'b0; 
    assign out[7692] = 1'b0; 
    assign out[7693] = 1'b0; 
    assign out[7694] = 1'b0; 
    assign out[7695] = 1'b0; 
    assign out[7696] = 1'b0; 
    assign out[7697] = 1'b0; 
    assign out[7698] = 1'b0; 
    assign out[7699] = 1'b0; 
    assign out[7700] = 1'b0; 
    assign out[7701] = 1'b0; 
    assign out[7702] = 1'b0; 
    assign out[7703] = 1'b0; 
    assign out[7704] = 1'b0; 
    assign out[7705] = 1'b0; 
    assign out[7706] = 1'b0; 
    assign out[7707] = 1'b0; 
    assign out[7708] = 1'b0; 
    assign out[7709] = 1'b0; 
    assign out[7710] = 1'b0; 
    assign out[7711] = 1'b0; 
    assign out[7712] = 1'b0; 
    assign out[7713] = 1'b0; 
    assign out[7714] = 1'b0; 
    assign out[7715] = 1'b0; 
    assign out[7716] = 1'b0; 
    assign out[7717] = 1'b0; 
    assign out[7718] = 1'b0; 
    assign out[7719] = 1'b0; 
    assign out[7720] = 1'b0; 
    assign out[7721] = 1'b0; 
    assign out[7722] = 1'b0; 
    assign out[7723] = 1'b0; 
    assign out[7724] = 1'b0; 
    assign out[7725] = 1'b0; 
    assign out[7726] = 1'b0; 
    assign out[7727] = 1'b0; 
    assign out[7728] = 1'b0; 
    assign out[7729] = 1'b0; 
    assign out[7730] = 1'b0; 
    assign out[7731] = 1'b0; 
    assign out[7732] = 1'b0; 
    assign out[7733] = 1'b0; 
    assign out[7734] = 1'b0; 
    assign out[7735] = 1'b0; 
    assign out[7736] = 1'b0; 
    assign out[7737] = 1'b0; 
    assign out[7738] = 1'b0; 
    assign out[7739] = 1'b0; 
    assign out[7740] = 1'b0; 
    assign out[7741] = 1'b0; 
    assign out[7742] = 1'b0; 
    assign out[7743] = 1'b0; 
    assign out[7744] = 1'b0; 
    assign out[7745] = 1'b0; 
    assign out[7746] = 1'b0; 
    assign out[7747] = 1'b0; 
    assign out[7748] = 1'b0; 
    assign out[7749] = 1'b0; 
    assign out[7750] = 1'b0; 
    assign out[7751] = 1'b0; 
    assign out[7752] = 1'b0; 
    assign out[7753] = 1'b0; 
    assign out[7754] = 1'b0; 
    assign out[7755] = 1'b0; 
    assign out[7756] = 1'b0; 
    assign out[7757] = 1'b0; 
    assign out[7758] = 1'b0; 
    assign out[7759] = 1'b0; 
    assign out[7760] = 1'b0; 
    assign out[7761] = 1'b0; 
    assign out[7762] = 1'b0; 
    assign out[7763] = 1'b0; 
    assign out[7764] = 1'b0; 
    assign out[7765] = 1'b0; 
    assign out[7766] = 1'b0; 
    assign out[7767] = 1'b0; 
    assign out[7768] = 1'b0; 
    assign out[7769] = 1'b0; 
    assign out[7770] = 1'b0; 
    assign out[7771] = 1'b0; 
    assign out[7772] = 1'b0; 
    assign out[7773] = 1'b0; 
    assign out[7774] = 1'b0; 
    assign out[7775] = 1'b0; 
    assign out[7776] = 1'b0; 
    assign out[7777] = 1'b0; 
    assign out[7778] = 1'b0; 
    assign out[7779] = 1'b0; 
    assign out[7780] = 1'b0; 
    assign out[7781] = 1'b0; 
    assign out[7782] = 1'b0; 
    assign out[7783] = 1'b0; 
    assign out[7784] = 1'b0; 
    assign out[7785] = 1'b0; 
    assign out[7786] = 1'b0; 
    assign out[7787] = 1'b0; 
    assign out[7788] = 1'b0; 
    assign out[7789] = 1'b0; 
    assign out[7790] = 1'b0; 
    assign out[7791] = 1'b0; 
    assign out[7792] = 1'b0; 
    assign out[7793] = 1'b0; 
    assign out[7794] = 1'b0; 
    assign out[7795] = 1'b0; 
    assign out[7796] = 1'b0; 
    assign out[7797] = 1'b0; 
    assign out[7798] = 1'b0; 
    assign out[7799] = 1'b0; 
    assign out[7800] = 1'b0; 
    assign out[7801] = 1'b0; 
    assign out[7802] = 1'b0; 
    assign out[7803] = 1'b0; 
    assign out[7804] = 1'b0; 
    assign out[7805] = 1'b0; 
    assign out[7806] = 1'b0; 
    assign out[7807] = 1'b0; 
    assign out[7808] = 1'b0; 
    assign out[7809] = 1'b0; 
    assign out[7810] = 1'b0; 
    assign out[7811] = 1'b0; 
    assign out[7812] = 1'b0; 
    assign out[7813] = 1'b0; 
    assign out[7814] = 1'b0; 
    assign out[7815] = 1'b0; 
    assign out[7816] = 1'b0; 
    assign out[7817] = 1'b0; 
    assign out[7818] = 1'b0; 
    assign out[7819] = 1'b0; 
    assign out[7820] = 1'b0; 
    assign out[7821] = 1'b0; 
    assign out[7822] = 1'b0; 
    assign out[7823] = 1'b0; 
    assign out[7824] = 1'b0; 
    assign out[7825] = 1'b0; 
    assign out[7826] = 1'b0; 
    assign out[7827] = 1'b0; 
    assign out[7828] = 1'b0; 
    assign out[7829] = 1'b0; 
    assign out[7830] = 1'b0; 
    assign out[7831] = 1'b0; 
    assign out[7832] = 1'b0; 
    assign out[7833] = 1'b0; 
    assign out[7834] = 1'b0; 
    assign out[7835] = 1'b0; 
    assign out[7836] = 1'b0; 
    assign out[7837] = 1'b0; 
    assign out[7838] = 1'b0; 
    assign out[7839] = 1'b0; 
    assign out[7840] = 1'b0; 
    assign out[7841] = 1'b0; 
    assign out[7842] = 1'b0; 
    assign out[7843] = 1'b0; 
    assign out[7844] = 1'b0; 
    assign out[7845] = 1'b0; 
    assign out[7846] = 1'b0; 
    assign out[7847] = 1'b0; 
    assign out[7848] = 1'b0; 
    assign out[7849] = 1'b0; 
    assign out[7850] = 1'b0; 
    assign out[7851] = 1'b0; 
    assign out[7852] = 1'b0; 
    assign out[7853] = 1'b0; 
    assign out[7854] = 1'b0; 
    assign out[7855] = 1'b0; 
    assign out[7856] = 1'b0; 
    assign out[7857] = 1'b0; 
    assign out[7858] = 1'b0; 
    assign out[7859] = 1'b0; 
    assign out[7860] = 1'b0; 
    assign out[7861] = 1'b0; 
    assign out[7862] = 1'b0; 
    assign out[7863] = 1'b0; 
    assign out[7864] = 1'b0; 
    assign out[7865] = 1'b0; 
    assign out[7866] = 1'b0; 
    assign out[7867] = 1'b0; 
    assign out[7868] = 1'b0; 
    assign out[7869] = 1'b0; 
    assign out[7870] = 1'b0; 
    assign out[7871] = 1'b0; 
    assign out[7872] = 1'b0; 
    assign out[7873] = 1'b0; 
    assign out[7874] = 1'b0; 
    assign out[7875] = 1'b0; 
    assign out[7876] = 1'b0; 
    assign out[7877] = 1'b0; 
    assign out[7878] = 1'b0; 
    assign out[7879] = 1'b0; 
    assign out[7880] = 1'b0; 
    assign out[7881] = 1'b0; 
    assign out[7882] = 1'b0; 
    assign out[7883] = 1'b0; 
    assign out[7884] = 1'b0; 
    assign out[7885] = 1'b0; 
    assign out[7886] = 1'b0; 
    assign out[7887] = 1'b0; 
    assign out[7888] = 1'b0; 
    assign out[7889] = 1'b0; 
    assign out[7890] = 1'b0; 
    assign out[7891] = 1'b0; 
    assign out[7892] = 1'b0; 
    assign out[7893] = 1'b0; 
    assign out[7894] = 1'b0; 
    assign out[7895] = 1'b0; 
    assign out[7896] = 1'b0; 
    assign out[7897] = 1'b0; 
    assign out[7898] = 1'b0; 
    assign out[7899] = 1'b0; 
    assign out[7900] = 1'b0; 
    assign out[7901] = 1'b0; 
    assign out[7902] = 1'b0; 
    assign out[7903] = 1'b0; 
    assign out[7904] = 1'b0; 
    assign out[7905] = 1'b0; 
    assign out[7906] = 1'b0; 
    assign out[7907] = 1'b0; 
    assign out[7908] = 1'b0; 
    assign out[7909] = 1'b0; 
    assign out[7910] = 1'b0; 
    assign out[7911] = 1'b0; 
    assign out[7912] = 1'b0; 
    assign out[7913] = 1'b0; 
    assign out[7914] = 1'b0; 
    assign out[7915] = 1'b0; 
    assign out[7916] = 1'b0; 
    assign out[7917] = 1'b0; 
    assign out[7918] = 1'b0; 
    assign out[7919] = 1'b0; 
    assign out[7920] = 1'b0; 
    assign out[7921] = 1'b0; 
    assign out[7922] = 1'b0; 
    assign out[7923] = 1'b0; 
    assign out[7924] = 1'b0; 
    assign out[7925] = 1'b0; 
    assign out[7926] = 1'b0; 
    assign out[7927] = 1'b0; 
    assign out[7928] = 1'b0; 
    assign out[7929] = 1'b0; 
    assign out[7930] = 1'b0; 
    assign out[7931] = 1'b0; 
    assign out[7932] = 1'b0; 
    assign out[7933] = 1'b0; 
    assign out[7934] = 1'b0; 
    assign out[7935] = 1'b0; 
    assign out[7936] = 1'b0; 
    assign out[7937] = 1'b0; 
    assign out[7938] = 1'b0; 
    assign out[7939] = 1'b0; 
    assign out[7940] = 1'b0; 
    assign out[7941] = 1'b0; 
    assign out[7942] = 1'b0; 
    assign out[7943] = 1'b0; 
    assign out[7944] = 1'b0; 
    assign out[7945] = 1'b0; 
    assign out[7946] = 1'b0; 
    assign out[7947] = 1'b0; 
    assign out[7948] = 1'b0; 
    assign out[7949] = 1'b0; 
    assign out[7950] = 1'b0; 
    assign out[7951] = 1'b0; 
    assign out[7952] = 1'b0; 
    assign out[7953] = 1'b0; 
    assign out[7954] = 1'b0; 
    assign out[7955] = 1'b0; 
    assign out[7956] = 1'b0; 
    assign out[7957] = 1'b0; 
    assign out[7958] = 1'b0; 
    assign out[7959] = 1'b0; 
    assign out[7960] = 1'b0; 
    assign out[7961] = 1'b0; 
    assign out[7962] = 1'b0; 
    assign out[7963] = 1'b0; 
    assign out[7964] = 1'b0; 
    assign out[7965] = 1'b0; 
    assign out[7966] = 1'b0; 
    assign out[7967] = 1'b0; 
    assign out[7968] = 1'b0; 
    assign out[7969] = 1'b0; 
    assign out[7970] = 1'b0; 
    assign out[7971] = 1'b0; 
    assign out[7972] = 1'b0; 
    assign out[7973] = 1'b0; 
    assign out[7974] = 1'b0; 
    assign out[7975] = 1'b0; 
    assign out[7976] = 1'b0; 
    assign out[7977] = 1'b0; 
    assign out[7978] = 1'b0; 
    assign out[7979] = 1'b0; 
    assign out[7980] = 1'b0; 
    assign out[7981] = 1'b0; 
    assign out[7982] = 1'b0; 
    assign out[7983] = 1'b0; 
    assign out[7984] = 1'b0; 
    assign out[7985] = 1'b0; 
    assign out[7986] = 1'b0; 
    assign out[7987] = 1'b0; 
    assign out[7988] = 1'b0; 
    assign out[7989] = 1'b0; 
    assign out[7990] = 1'b0; 
    assign out[7991] = 1'b0; 
    assign out[7992] = 1'b0; 
    assign out[7993] = 1'b0; 
    assign out[7994] = 1'b0; 
    assign out[7995] = 1'b0; 
    assign out[7996] = 1'b0; 
    assign out[7997] = 1'b0; 
    assign out[7998] = 1'b0; 
    assign out[7999] = 1'b0; 
    // Arrange outputs in categories ================================================
    assign categories[5109:0] = out[5109:0];

endmodule
