// Generated from: 20251204-084921_binTestAcc8873_seed190838_epochs100_2x12000_b256_lr50_interconnect.npz

module net (
    input  wire [1023:0] in,
    output wire [11999:0] out,
    output wire [7999:0] categories
);
    wire [11999:0] layer_0;

    // Layer 0 ============================================================
    assign layer_0[0] = in[502] & in[186]; 
    assign layer_0[1] = in[872]; 
    assign layer_0[2] = in[596] | in[830]; 
    assign layer_0[3] = ~(in[713] ^ in[835]); 
    assign layer_0[4] = in[164] & ~in[162]; 
    assign layer_0[5] = ~(in[577] ^ in[469]); 
    assign layer_0[6] = in[435] ^ in[793]; 
    assign layer_0[7] = ~(in[843] & in[11]); 
    assign layer_0[8] = in[551] ^ in[300]; 
    assign layer_0[9] = ~(in[342] ^ in[845]); 
    assign layer_0[10] = in[970] ^ in[512]; 
    assign layer_0[11] = ~(in[18] | in[738]); 
    assign layer_0[12] = ~(in[284] | in[683]); 
    assign layer_0[13] = ~(in[963] | in[549]); 
    assign layer_0[14] = in[443] & in[100]; 
    assign layer_0[15] = in[145] & in[73]; 
    assign layer_0[16] = ~in[892]; 
    assign layer_0[17] = in[21]; 
    assign layer_0[18] = in[84] & ~in[473]; 
    assign layer_0[19] = ~in[354] | (in[797] & in[354]); 
    assign layer_0[20] = in[985] ^ in[595]; 
    assign layer_0[21] = ~(in[110] ^ in[74]); 
    assign layer_0[22] = 1'b0; 
    assign layer_0[23] = ~in[936]; 
    assign layer_0[24] = ~in[229] | (in[461] & in[229]); 
    assign layer_0[25] = 1'b0; 
    assign layer_0[26] = ~(in[570] & in[183]); 
    assign layer_0[27] = in[483]; 
    assign layer_0[28] = ~(in[193] & in[192]); 
    assign layer_0[29] = in[419] & ~in[55]; 
    assign layer_0[30] = in[697] & ~in[862]; 
    assign layer_0[31] = in[84] & ~in[604]; 
    assign layer_0[32] = ~(in[595] & in[368]); 
    assign layer_0[33] = ~in[709]; 
    assign layer_0[34] = ~(in[760] ^ in[758]); 
    assign layer_0[35] = in[666] & in[346]; 
    assign layer_0[36] = in[338] ^ in[292]; 
    assign layer_0[37] = ~in[207]; 
    assign layer_0[38] = ~in[533] | (in[638] & in[533]); 
    assign layer_0[39] = ~in[484]; 
    assign layer_0[40] = in[85] & ~in[1007]; 
    assign layer_0[41] = ~in[552] | (in[554] & in[552]); 
    assign layer_0[42] = in[872] & in[920]; 
    assign layer_0[43] = in[516]; 
    assign layer_0[44] = in[601] & in[456]; 
    assign layer_0[45] = ~(in[630] & in[621]); 
    assign layer_0[46] = in[244]; 
    assign layer_0[47] = ~in[967] | (in[940] & in[967]); 
    assign layer_0[48] = in[823] ^ in[20]; 
    assign layer_0[49] = ~in[203]; 
    assign layer_0[50] = in[919] & ~in[957]; 
    assign layer_0[51] = ~in[276]; 
    assign layer_0[52] = ~(in[828] ^ in[940]); 
    assign layer_0[53] = in[889] & ~in[728]; 
    assign layer_0[54] = in[102] & ~in[121]; 
    assign layer_0[55] = in[745] ^ in[194]; 
    assign layer_0[56] = ~(in[271] | in[141]); 
    assign layer_0[57] = ~in[316] | (in[316] & in[975]); 
    assign layer_0[58] = ~(in[656] ^ in[670]); 
    assign layer_0[59] = ~(in[110] ^ in[885]); 
    assign layer_0[60] = in[956]; 
    assign layer_0[61] = in[502]; 
    assign layer_0[62] = ~in[421] | (in[55] & in[421]); 
    assign layer_0[63] = ~(in[1017] ^ in[147]); 
    assign layer_0[64] = in[488] & ~in[541]; 
    assign layer_0[65] = in[1008] | in[233]; 
    assign layer_0[66] = in[551] & ~in[779]; 
    assign layer_0[67] = ~in[239]; 
    assign layer_0[68] = in[787]; 
    assign layer_0[69] = ~in[98] | (in[98] & in[96]); 
    assign layer_0[70] = in[397] ^ in[386]; 
    assign layer_0[71] = ~in[50] | (in[490] & in[50]); 
    assign layer_0[72] = ~(in[67] ^ in[709]); 
    assign layer_0[73] = in[440]; 
    assign layer_0[74] = ~in[342]; 
    assign layer_0[75] = in[475]; 
    assign layer_0[76] = in[775] & in[75]; 
    assign layer_0[77] = in[597] & ~in[835]; 
    assign layer_0[78] = in[738] & ~in[490]; 
    assign layer_0[79] = in[343]; 
    assign layer_0[80] = in[332] ^ in[970]; 
    assign layer_0[81] = in[104] & ~in[462]; 
    assign layer_0[82] = in[471] ^ in[689]; 
    assign layer_0[83] = ~(in[712] ^ in[713]); 
    assign layer_0[84] = in[649]; 
    assign layer_0[85] = in[791] | in[1011]; 
    assign layer_0[86] = in[282] & in[3]; 
    assign layer_0[87] = ~(in[701] | in[603]); 
    assign layer_0[88] = ~(in[403] & in[102]); 
    assign layer_0[89] = in[78]; 
    assign layer_0[90] = ~(in[307] | in[66]); 
    assign layer_0[91] = ~(in[278] & in[661]); 
    assign layer_0[92] = ~(in[518] ^ in[520]); 
    assign layer_0[93] = ~(in[14] ^ in[917]); 
    assign layer_0[94] = ~(in[28] ^ in[652]); 
    assign layer_0[95] = ~(in[192] ^ in[755]); 
    assign layer_0[96] = ~(in[494] ^ in[907]); 
    assign layer_0[97] = in[920] & ~in[823]; 
    assign layer_0[98] = ~(in[870] ^ in[792]); 
    assign layer_0[99] = in[888] ^ in[906]; 
    assign layer_0[100] = ~in[428]; 
    assign layer_0[101] = ~(in[2] ^ in[283]); 
    assign layer_0[102] = in[534] & in[475]; 
    assign layer_0[103] = in[692] & ~in[743]; 
    assign layer_0[104] = in[294]; 
    assign layer_0[105] = ~(in[111] ^ in[556]); 
    assign layer_0[106] = ~(in[587] | in[99]); 
    assign layer_0[107] = in[501] & in[388]; 
    assign layer_0[108] = ~(in[769] ^ in[448]); 
    assign layer_0[109] = ~(in[627] ^ in[165]); 
    assign layer_0[110] = in[92] & ~in[981]; 
    assign layer_0[111] = ~in[988] | (in[330] & in[988]); 
    assign layer_0[112] = ~in[910] | (in[947] & in[910]); 
    assign layer_0[113] = in[346] & ~in[533]; 
    assign layer_0[114] = ~in[78]; 
    assign layer_0[115] = in[740] ^ in[599]; 
    assign layer_0[116] = in[618]; 
    assign layer_0[117] = in[731]; 
    assign layer_0[118] = ~(in[891] ^ in[459]); 
    assign layer_0[119] = in[416] ^ in[952]; 
    assign layer_0[120] = ~in[623]; 
    assign layer_0[121] = ~(in[96] ^ in[205]); 
    assign layer_0[122] = in[629] ^ in[875]; 
    assign layer_0[123] = in[729]; 
    assign layer_0[124] = in[156]; 
    assign layer_0[125] = 1'b1; 
    assign layer_0[126] = ~(in[275] ^ in[237]); 
    assign layer_0[127] = in[194] ^ in[570]; 
    assign layer_0[128] = in[347] & in[580]; 
    assign layer_0[129] = in[427]; 
    assign layer_0[130] = ~in[424]; 
    assign layer_0[131] = in[1003]; 
    assign layer_0[132] = in[509] ^ in[318]; 
    assign layer_0[133] = ~(in[537] | in[577]); 
    assign layer_0[134] = in[38]; 
    assign layer_0[135] = ~(in[894] & in[861]); 
    assign layer_0[136] = in[532] & in[210]; 
    assign layer_0[137] = ~in[878] | (in[878] & in[984]); 
    assign layer_0[138] = 1'b1; 
    assign layer_0[139] = ~in[12]; 
    assign layer_0[140] = in[220] & ~in[723]; 
    assign layer_0[141] = ~(in[52] & in[537]); 
    assign layer_0[142] = ~(in[613] ^ in[68]); 
    assign layer_0[143] = in[409] | in[1019]; 
    assign layer_0[144] = ~in[836]; 
    assign layer_0[145] = in[730]; 
    assign layer_0[146] = 1'b0; 
    assign layer_0[147] = ~(in[275] ^ in[714]); 
    assign layer_0[148] = ~in[463] | (in[260] & in[463]); 
    assign layer_0[149] = ~in[622]; 
    assign layer_0[150] = in[725]; 
    assign layer_0[151] = ~in[38]; 
    assign layer_0[152] = ~(in[549] ^ in[493]); 
    assign layer_0[153] = in[900] & ~in[897]; 
    assign layer_0[154] = in[485] ^ in[939]; 
    assign layer_0[155] = ~in[855] | (in[855] & in[891]); 
    assign layer_0[156] = ~(in[999] ^ in[173]); 
    assign layer_0[157] = in[74]; 
    assign layer_0[158] = in[906] ^ in[187]; 
    assign layer_0[159] = ~(in[996] ^ in[506]); 
    assign layer_0[160] = ~(in[934] ^ in[680]); 
    assign layer_0[161] = ~in[107] | (in[107] & in[92]); 
    assign layer_0[162] = in[695]; 
    assign layer_0[163] = ~(in[365] ^ in[45]); 
    assign layer_0[164] = ~in[395] | (in[395] & in[123]); 
    assign layer_0[165] = in[295] & ~in[755]; 
    assign layer_0[166] = in[910]; 
    assign layer_0[167] = ~(in[24] ^ in[764]); 
    assign layer_0[168] = 1'b1; 
    assign layer_0[169] = ~(in[361] ^ in[875]); 
    assign layer_0[170] = ~(in[461] ^ in[598]); 
    assign layer_0[171] = in[565] & ~in[777]; 
    assign layer_0[172] = ~in[489] | (in[489] & in[840]); 
    assign layer_0[173] = in[29] | in[464]; 
    assign layer_0[174] = ~(in[806] ^ in[459]); 
    assign layer_0[175] = in[550] ^ in[520]; 
    assign layer_0[176] = in[966] ^ in[904]; 
    assign layer_0[177] = in[633]; 
    assign layer_0[178] = 1'b1; 
    assign layer_0[179] = in[726] & ~in[783]; 
    assign layer_0[180] = in[397] & in[915]; 
    assign layer_0[181] = in[23] & in[412]; 
    assign layer_0[182] = ~(in[90] ^ in[587]); 
    assign layer_0[183] = ~(in[681] ^ in[941]); 
    assign layer_0[184] = in[1018] | in[912]; 
    assign layer_0[185] = in[317]; 
    assign layer_0[186] = in[59] & ~in[177]; 
    assign layer_0[187] = in[507]; 
    assign layer_0[188] = ~(in[963] ^ in[597]); 
    assign layer_0[189] = 1'b0; 
    assign layer_0[190] = in[599] & ~in[740]; 
    assign layer_0[191] = ~(in[553] ^ in[76]); 
    assign layer_0[192] = ~(in[483] ^ in[140]); 
    assign layer_0[193] = in[840] | in[952]; 
    assign layer_0[194] = in[952]; 
    assign layer_0[195] = in[474] & ~in[603]; 
    assign layer_0[196] = in[903] | in[605]; 
    assign layer_0[197] = in[748] & ~in[408]; 
    assign layer_0[198] = in[570] & ~in[371]; 
    assign layer_0[199] = in[21]; 
    assign layer_0[200] = in[593] | in[114]; 
    assign layer_0[201] = ~(in[654] ^ in[172]); 
    assign layer_0[202] = ~in[581]; 
    assign layer_0[203] = in[722] ^ in[673]; 
    assign layer_0[204] = ~in[419] | (in[37] & in[419]); 
    assign layer_0[205] = in[457] & in[506]; 
    assign layer_0[206] = in[506] & ~in[13]; 
    assign layer_0[207] = ~in[877] | (in[877] & in[726]); 
    assign layer_0[208] = ~(in[950] ^ in[968]); 
    assign layer_0[209] = ~(in[677] ^ in[222]); 
    assign layer_0[210] = in[109] & ~in[154]; 
    assign layer_0[211] = ~(in[612] ^ in[603]); 
    assign layer_0[212] = ~(in[1004] | in[871]); 
    assign layer_0[213] = in[483] & in[508]; 
    assign layer_0[214] = in[475]; 
    assign layer_0[215] = in[684] & in[339]; 
    assign layer_0[216] = ~in[279] | (in[279] & in[19]); 
    assign layer_0[217] = ~(in[745] ^ in[647]); 
    assign layer_0[218] = in[660]; 
    assign layer_0[219] = in[498]; 
    assign layer_0[220] = ~(in[82] & in[88]); 
    assign layer_0[221] = ~(in[65] ^ in[1002]); 
    assign layer_0[222] = in[375] & ~in[772]; 
    assign layer_0[223] = ~(in[440] | in[688]); 
    assign layer_0[224] = ~in[193]; 
    assign layer_0[225] = ~(in[154] & in[488]); 
    assign layer_0[226] = in[980] ^ in[70]; 
    assign layer_0[227] = in[115]; 
    assign layer_0[228] = in[210] & ~in[18]; 
    assign layer_0[229] = in[950] ^ in[579]; 
    assign layer_0[230] = ~(in[966] ^ in[986]); 
    assign layer_0[231] = in[886] ^ in[55]; 
    assign layer_0[232] = in[209] & in[613]; 
    assign layer_0[233] = ~(in[62] & in[549]); 
    assign layer_0[234] = ~in[580]; 
    assign layer_0[235] = in[206] ^ in[15]; 
    assign layer_0[236] = in[238] ^ in[262]; 
    assign layer_0[237] = in[473] ^ in[784]; 
    assign layer_0[238] = ~(in[1002] ^ in[52]); 
    assign layer_0[239] = ~(in[936] ^ in[444]); 
    assign layer_0[240] = in[534]; 
    assign layer_0[241] = ~(in[882] & in[964]); 
    assign layer_0[242] = in[904] | in[232]; 
    assign layer_0[243] = ~(in[506] ^ in[871]); 
    assign layer_0[244] = ~(in[838] ^ in[550]); 
    assign layer_0[245] = ~(in[466] | in[991]); 
    assign layer_0[246] = ~in[611]; 
    assign layer_0[247] = ~in[280]; 
    assign layer_0[248] = in[139] & ~in[482]; 
    assign layer_0[249] = ~(in[753] | in[342]); 
    assign layer_0[250] = 1'b1; 
    assign layer_0[251] = in[257]; 
    assign layer_0[252] = ~(in[35] | in[544]); 
    assign layer_0[253] = in[564] & ~in[618]; 
    assign layer_0[254] = 1'b0; 
    assign layer_0[255] = in[909] ^ in[97]; 
    assign layer_0[256] = ~(in[273] ^ in[1015]); 
    assign layer_0[257] = ~(in[115] | in[944]); 
    assign layer_0[258] = ~(in[650] ^ in[679]); 
    assign layer_0[259] = ~(in[924] ^ in[993]); 
    assign layer_0[260] = ~in[508]; 
    assign layer_0[261] = in[590] ^ in[462]; 
    assign layer_0[262] = in[894] & ~in[719]; 
    assign layer_0[263] = in[668]; 
    assign layer_0[264] = in[110]; 
    assign layer_0[265] = in[703] & in[87]; 
    assign layer_0[266] = in[123] ^ in[349]; 
    assign layer_0[267] = in[696] & in[944]; 
    assign layer_0[268] = in[240] & ~in[871]; 
    assign layer_0[269] = ~in[936] | (in[415] & in[936]); 
    assign layer_0[270] = 1'b1; 
    assign layer_0[271] = in[75] ^ in[612]; 
    assign layer_0[272] = in[629] ^ in[883]; 
    assign layer_0[273] = in[265] | in[283]; 
    assign layer_0[274] = ~(in[940] ^ in[29]); 
    assign layer_0[275] = in[724] ^ in[905]; 
    assign layer_0[276] = in[548] & in[542]; 
    assign layer_0[277] = in[709]; 
    assign layer_0[278] = in[649] | in[991]; 
    assign layer_0[279] = ~in[858] | (in[637] & in[858]); 
    assign layer_0[280] = in[32]; 
    assign layer_0[281] = ~(in[716] ^ in[505]); 
    assign layer_0[282] = ~in[844] | (in[844] & in[930]); 
    assign layer_0[283] = in[371] | in[947]; 
    assign layer_0[284] = ~(in[920] ^ in[571]); 
    assign layer_0[285] = ~in[260]; 
    assign layer_0[286] = ~in[413]; 
    assign layer_0[287] = ~(in[30] | in[306]); 
    assign layer_0[288] = ~(in[488] & in[82]); 
    assign layer_0[289] = ~(in[860] & in[926]); 
    assign layer_0[290] = in[101] ^ in[75]; 
    assign layer_0[291] = in[203] & ~in[357]; 
    assign layer_0[292] = ~(in[934] | in[231]); 
    assign layer_0[293] = ~(in[621] ^ in[690]); 
    assign layer_0[294] = in[742] ^ in[898]; 
    assign layer_0[295] = in[328] & ~in[550]; 
    assign layer_0[296] = ~(in[790] ^ in[964]); 
    assign layer_0[297] = ~in[113]; 
    assign layer_0[298] = in[195]; 
    assign layer_0[299] = in[517] | in[531]; 
    assign layer_0[300] = in[6] & ~in[143]; 
    assign layer_0[301] = in[5] ^ in[229]; 
    assign layer_0[302] = in[160] & ~in[982]; 
    assign layer_0[303] = in[647]; 
    assign layer_0[304] = ~(in[463] ^ in[606]); 
    assign layer_0[305] = ~in[649] | (in[649] & in[900]); 
    assign layer_0[306] = ~(in[1002] ^ in[42]); 
    assign layer_0[307] = in[2] ^ in[470]; 
    assign layer_0[308] = ~(in[757] ^ in[661]); 
    assign layer_0[309] = in[297] ^ in[222]; 
    assign layer_0[310] = ~(in[1001] | in[242]); 
    assign layer_0[311] = ~(in[860] ^ in[849]); 
    assign layer_0[312] = in[844] ^ in[37]; 
    assign layer_0[313] = in[243]; 
    assign layer_0[314] = ~(in[374] & in[51]); 
    assign layer_0[315] = ~in[656] | (in[500] & in[656]); 
    assign layer_0[316] = in[634] ^ in[648]; 
    assign layer_0[317] = ~(in[725] ^ in[873]); 
    assign layer_0[318] = ~in[862]; 
    assign layer_0[319] = ~(in[968] ^ in[872]); 
    assign layer_0[320] = in[856] ^ in[478]; 
    assign layer_0[321] = ~in[951] | (in[450] & in[951]); 
    assign layer_0[322] = in[724] ^ in[599]; 
    assign layer_0[323] = in[893] & ~in[584]; 
    assign layer_0[324] = ~in[472]; 
    assign layer_0[325] = in[704] ^ in[967]; 
    assign layer_0[326] = in[334] & ~in[851]; 
    assign layer_0[327] = in[292] & ~in[1010]; 
    assign layer_0[328] = ~(in[157] | in[875]); 
    assign layer_0[329] = in[809] & ~in[788]; 
    assign layer_0[330] = ~in[664] | (in[664] & in[1017]); 
    assign layer_0[331] = in[943]; 
    assign layer_0[332] = ~(in[631] | in[300]); 
    assign layer_0[333] = ~in[740] | (in[740] & in[976]); 
    assign layer_0[334] = ~(in[113] & in[58]); 
    assign layer_0[335] = ~in[373] | (in[350] & in[373]); 
    assign layer_0[336] = ~in[115] | (in[115] & in[349]); 
    assign layer_0[337] = ~(in[929] ^ in[463]); 
    assign layer_0[338] = ~(in[987] ^ in[956]); 
    assign layer_0[339] = ~(in[700] | in[147]); 
    assign layer_0[340] = in[813]; 
    assign layer_0[341] = in[770] ^ in[791]; 
    assign layer_0[342] = in[447] & in[436]; 
    assign layer_0[343] = ~(in[267] ^ in[981]); 
    assign layer_0[344] = in[714] ^ in[504]; 
    assign layer_0[345] = ~(in[354] ^ in[973]); 
    assign layer_0[346] = in[760] ^ in[507]; 
    assign layer_0[347] = ~in[202]; 
    assign layer_0[348] = in[506] | in[949]; 
    assign layer_0[349] = ~(in[205] & in[622]); 
    assign layer_0[350] = in[924]; 
    assign layer_0[351] = ~in[958] | (in[958] & in[607]); 
    assign layer_0[352] = ~(in[95] ^ in[309]); 
    assign layer_0[353] = ~in[861]; 
    assign layer_0[354] = ~(in[921] ^ in[824]); 
    assign layer_0[355] = in[622] ^ in[853]; 
    assign layer_0[356] = ~in[77] | (in[77] & in[460]); 
    assign layer_0[357] = ~in[922] | (in[922] & in[845]); 
    assign layer_0[358] = ~in[423]; 
    assign layer_0[359] = in[387]; 
    assign layer_0[360] = in[631] ^ in[600]; 
    assign layer_0[361] = ~(in[354] | in[553]); 
    assign layer_0[362] = in[172] ^ in[285]; 
    assign layer_0[363] = in[778] ^ in[13]; 
    assign layer_0[364] = ~(in[451] ^ in[966]); 
    assign layer_0[365] = in[715] & ~in[596]; 
    assign layer_0[366] = ~(in[277] ^ in[493]); 
    assign layer_0[367] = ~(in[790] ^ in[806]); 
    assign layer_0[368] = ~(in[322] ^ in[607]); 
    assign layer_0[369] = in[794]; 
    assign layer_0[370] = ~in[1013] | (in[1013] & in[301]); 
    assign layer_0[371] = ~(in[586] ^ in[890]); 
    assign layer_0[372] = ~(in[483] & in[152]); 
    assign layer_0[373] = ~(in[863] ^ in[349]); 
    assign layer_0[374] = in[507] ^ in[92]; 
    assign layer_0[375] = in[631] ^ in[729]; 
    assign layer_0[376] = 1'b0; 
    assign layer_0[377] = in[556] & ~in[947]; 
    assign layer_0[378] = ~in[400] | (in[400] & in[800]); 
    assign layer_0[379] = ~(in[952] ^ in[954]); 
    assign layer_0[380] = in[218]; 
    assign layer_0[381] = in[477] ^ in[333]; 
    assign layer_0[382] = in[583] | in[610]; 
    assign layer_0[383] = ~(in[936] ^ in[937]); 
    assign layer_0[384] = ~in[598] | (in[598] & in[572]); 
    assign layer_0[385] = in[220]; 
    assign layer_0[386] = ~(in[938] ^ in[922]); 
    assign layer_0[387] = ~in[500] | (in[356] & in[500]); 
    assign layer_0[388] = ~(in[697] ^ in[505]); 
    assign layer_0[389] = in[892] & ~in[111]; 
    assign layer_0[390] = in[252]; 
    assign layer_0[391] = in[1] | in[683]; 
    assign layer_0[392] = in[395]; 
    assign layer_0[393] = in[174] | in[523]; 
    assign layer_0[394] = in[870]; 
    assign layer_0[395] = in[420]; 
    assign layer_0[396] = ~(in[966] | in[826]); 
    assign layer_0[397] = in[752] ^ in[540]; 
    assign layer_0[398] = ~(in[535] & in[584]); 
    assign layer_0[399] = ~(in[860] | in[859]); 
    assign layer_0[400] = in[857]; 
    assign layer_0[401] = ~in[975]; 
    assign layer_0[402] = in[933] ^ in[685]; 
    assign layer_0[403] = in[932] | in[1001]; 
    assign layer_0[404] = ~(in[268] ^ in[939]); 
    assign layer_0[405] = in[894] & ~in[611]; 
    assign layer_0[406] = ~in[700]; 
    assign layer_0[407] = ~(in[651] ^ in[268]); 
    assign layer_0[408] = ~(in[755] ^ in[995]); 
    assign layer_0[409] = ~(in[988] ^ in[857]); 
    assign layer_0[410] = in[332] ^ in[715]; 
    assign layer_0[411] = ~(in[761] ^ in[760]); 
    assign layer_0[412] = in[1016]; 
    assign layer_0[413] = ~(in[952] ^ in[904]); 
    assign layer_0[414] = in[272] | in[664]; 
    assign layer_0[415] = ~(in[902] ^ in[754]); 
    assign layer_0[416] = in[937] | in[10]; 
    assign layer_0[417] = in[585] | in[671]; 
    assign layer_0[418] = in[57] | in[816]; 
    assign layer_0[419] = in[866]; 
    assign layer_0[420] = in[312] & in[599]; 
    assign layer_0[421] = in[793] ^ in[873]; 
    assign layer_0[422] = ~(in[669] ^ in[207]); 
    assign layer_0[423] = in[634] & ~in[806]; 
    assign layer_0[424] = in[580] ^ in[444]; 
    assign layer_0[425] = ~in[217]; 
    assign layer_0[426] = ~(in[449] & in[751]); 
    assign layer_0[427] = ~(in[435] & in[428]); 
    assign layer_0[428] = in[904] ^ in[720]; 
    assign layer_0[429] = 1'b1; 
    assign layer_0[430] = ~(in[854] ^ in[240]); 
    assign layer_0[431] = in[599] & ~in[466]; 
    assign layer_0[432] = ~in[886]; 
    assign layer_0[433] = in[623]; 
    assign layer_0[434] = ~(in[848] ^ in[254]); 
    assign layer_0[435] = ~(in[1010] | in[657]); 
    assign layer_0[436] = ~(in[922] | in[238]); 
    assign layer_0[437] = ~(in[719] & in[143]); 
    assign layer_0[438] = in[954] | in[469]; 
    assign layer_0[439] = in[210] & in[189]; 
    assign layer_0[440] = ~(in[581] ^ in[1013]); 
    assign layer_0[441] = in[859] ^ in[500]; 
    assign layer_0[442] = in[715] & in[953]; 
    assign layer_0[443] = ~(in[409] & in[335]); 
    assign layer_0[444] = ~(in[450] ^ in[677]); 
    assign layer_0[445] = ~(in[964] ^ in[743]); 
    assign layer_0[446] = in[264] ^ in[981]; 
    assign layer_0[447] = ~(in[726] ^ in[65]); 
    assign layer_0[448] = ~in[566] | (in[508] & in[566]); 
    assign layer_0[449] = 1'b0; 
    assign layer_0[450] = ~in[264] | (in[264] & in[996]); 
    assign layer_0[451] = ~(in[147] & in[13]); 
    assign layer_0[452] = in[454] & in[77]; 
    assign layer_0[453] = in[888] & in[667]; 
    assign layer_0[454] = in[519] ^ in[549]; 
    assign layer_0[455] = ~in[854] | (in[854] & in[814]); 
    assign layer_0[456] = in[612] ^ in[855]; 
    assign layer_0[457] = ~in[254]; 
    assign layer_0[458] = in[236] & ~in[268]; 
    assign layer_0[459] = in[536] & ~in[797]; 
    assign layer_0[460] = ~(in[467] ^ in[301]); 
    assign layer_0[461] = in[841] ^ in[837]; 
    assign layer_0[462] = in[876]; 
    assign layer_0[463] = ~in[651] | (in[651] & in[576]); 
    assign layer_0[464] = in[642] ^ in[485]; 
    assign layer_0[465] = ~in[393] | (in[393] & in[937]); 
    assign layer_0[466] = in[534] | in[356]; 
    assign layer_0[467] = in[949] ^ in[57]; 
    assign layer_0[468] = in[840] & ~in[400]; 
    assign layer_0[469] = ~(in[520] | in[828]); 
    assign layer_0[470] = ~(in[443] ^ in[315]); 
    assign layer_0[471] = in[551] & ~in[306]; 
    assign layer_0[472] = ~(in[645] & in[538]); 
    assign layer_0[473] = ~in[300] | (in[300] & in[471]); 
    assign layer_0[474] = ~in[213]; 
    assign layer_0[475] = ~in[964] | (in[964] & in[871]); 
    assign layer_0[476] = ~(in[265] & in[730]); 
    assign layer_0[477] = in[936] ^ in[466]; 
    assign layer_0[478] = in[568] & ~in[773]; 
    assign layer_0[479] = ~in[23]; 
    assign layer_0[480] = ~in[173] | (in[635] & in[173]); 
    assign layer_0[481] = in[473] & ~in[84]; 
    assign layer_0[482] = in[385] & ~in[1022]; 
    assign layer_0[483] = in[201]; 
    assign layer_0[484] = ~(in[858] & in[923]); 
    assign layer_0[485] = in[601] & ~in[899]; 
    assign layer_0[486] = ~in[841]; 
    assign layer_0[487] = ~(in[912] ^ in[444]); 
    assign layer_0[488] = ~(in[55] ^ in[189]); 
    assign layer_0[489] = ~(in[43] ^ in[949]); 
    assign layer_0[490] = in[706]; 
    assign layer_0[491] = ~in[48] | (in[433] & in[48]); 
    assign layer_0[492] = ~(in[952] ^ in[371]); 
    assign layer_0[493] = ~(in[845] & in[359]); 
    assign layer_0[494] = in[517] ^ in[603]; 
    assign layer_0[495] = in[127] ^ in[891]; 
    assign layer_0[496] = in[445] | in[19]; 
    assign layer_0[497] = ~in[998] | (in[998] & in[781]); 
    assign layer_0[498] = in[669] | in[446]; 
    assign layer_0[499] = ~(in[429] ^ in[62]); 
    assign layer_0[500] = ~(in[471] & in[365]); 
    assign layer_0[501] = in[477] ^ in[469]; 
    assign layer_0[502] = in[212] & in[520]; 
    assign layer_0[503] = in[224]; 
    assign layer_0[504] = 1'b0; 
    assign layer_0[505] = in[244] ^ in[920]; 
    assign layer_0[506] = in[629]; 
    assign layer_0[507] = ~(in[963] ^ in[766]); 
    assign layer_0[508] = in[307] ^ in[882]; 
    assign layer_0[509] = in[623] & ~in[311]; 
    assign layer_0[510] = ~(in[657] ^ in[368]); 
    assign layer_0[511] = in[598]; 
    assign layer_0[512] = in[116] & in[618]; 
    assign layer_0[513] = in[29]; 
    assign layer_0[514] = in[983] & ~in[583]; 
    assign layer_0[515] = in[794] ^ in[99]; 
    assign layer_0[516] = ~(in[353] | in[831]); 
    assign layer_0[517] = ~in[615] | (in[485] & in[615]); 
    assign layer_0[518] = in[297]; 
    assign layer_0[519] = ~(in[4] | in[913]); 
    assign layer_0[520] = ~in[563] | (in[721] & in[563]); 
    assign layer_0[521] = ~in[436] | (in[160] & in[436]); 
    assign layer_0[522] = ~(in[918] | in[628]); 
    assign layer_0[523] = in[819] & ~in[343]; 
    assign layer_0[524] = in[599]; 
    assign layer_0[525] = ~(in[490] & in[739]); 
    assign layer_0[526] = in[775] ^ in[3]; 
    assign layer_0[527] = in[649] ^ in[638]; 
    assign layer_0[528] = in[856] ^ in[998]; 
    assign layer_0[529] = ~(in[900] & in[441]); 
    assign layer_0[530] = in[641] & ~in[557]; 
    assign layer_0[531] = ~(in[78] ^ in[222]); 
    assign layer_0[532] = in[906] & in[119]; 
    assign layer_0[533] = in[696]; 
    assign layer_0[534] = in[889] & ~in[13]; 
    assign layer_0[535] = ~(in[210] & in[236]); 
    assign layer_0[536] = in[62] ^ in[353]; 
    assign layer_0[537] = ~in[376]; 
    assign layer_0[538] = ~(in[839] | in[1018]); 
    assign layer_0[539] = in[932] ^ in[372]; 
    assign layer_0[540] = ~in[633]; 
    assign layer_0[541] = ~(in[716] ^ in[99]); 
    assign layer_0[542] = in[414] & ~in[649]; 
    assign layer_0[543] = in[314] & ~in[1002]; 
    assign layer_0[544] = ~in[205] | (in[760] & in[205]); 
    assign layer_0[545] = ~(in[168] & in[465]); 
    assign layer_0[546] = in[654]; 
    assign layer_0[547] = ~in[232] | (in[259] & in[232]); 
    assign layer_0[548] = in[807]; 
    assign layer_0[549] = in[639] | in[322]; 
    assign layer_0[550] = ~(in[824] ^ in[825]); 
    assign layer_0[551] = in[822] & ~in[591]; 
    assign layer_0[552] = in[16] ^ in[533]; 
    assign layer_0[553] = in[260] ^ in[937]; 
    assign layer_0[554] = ~(in[276] & in[573]); 
    assign layer_0[555] = ~(in[836] ^ in[276]); 
    assign layer_0[556] = in[355]; 
    assign layer_0[557] = in[438]; 
    assign layer_0[558] = in[952] ^ in[981]; 
    assign layer_0[559] = in[502] ^ in[733]; 
    assign layer_0[560] = ~(in[904] | in[887]); 
    assign layer_0[561] = ~(in[421] | in[873]); 
    assign layer_0[562] = ~(in[460] ^ in[660]); 
    assign layer_0[563] = ~(in[205] | in[758]); 
    assign layer_0[564] = ~(in[35] & in[438]); 
    assign layer_0[565] = in[704] ^ in[616]; 
    assign layer_0[566] = ~(in[587] ^ in[612]); 
    assign layer_0[567] = ~in[739] | (in[116] & in[739]); 
    assign layer_0[568] = ~in[689]; 
    assign layer_0[569] = ~(in[730] | in[309]); 
    assign layer_0[570] = ~(in[966] ^ in[968]); 
    assign layer_0[571] = in[481] ^ in[130]; 
    assign layer_0[572] = in[331] & in[67]; 
    assign layer_0[573] = in[613] & ~in[97]; 
    assign layer_0[574] = in[110]; 
    assign layer_0[575] = in[466] | in[791]; 
    assign layer_0[576] = ~(in[871] ^ in[873]); 
    assign layer_0[577] = ~(in[568] ^ in[931]); 
    assign layer_0[578] = in[824] ^ in[692]; 
    assign layer_0[579] = in[326] ^ in[590]; 
    assign layer_0[580] = ~in[942] | (in[880] & in[942]); 
    assign layer_0[581] = ~in[82]; 
    assign layer_0[582] = ~(in[1005] ^ in[723]); 
    assign layer_0[583] = in[95] & ~in[271]; 
    assign layer_0[584] = ~in[104]; 
    assign layer_0[585] = in[51] & ~in[306]; 
    assign layer_0[586] = ~in[620]; 
    assign layer_0[587] = ~(in[35] ^ in[968]); 
    assign layer_0[588] = in[355] | in[588]; 
    assign layer_0[589] = in[519] ^ in[619]; 
    assign layer_0[590] = in[699]; 
    assign layer_0[591] = in[204]; 
    assign layer_0[592] = ~(in[912] | in[704]); 
    assign layer_0[593] = in[901] ^ in[964]; 
    assign layer_0[594] = in[894] | in[933]; 
    assign layer_0[595] = in[680] & ~in[779]; 
    assign layer_0[596] = ~(in[972] & in[729]); 
    assign layer_0[597] = in[96] | in[553]; 
    assign layer_0[598] = ~(in[49] ^ in[909]); 
    assign layer_0[599] = ~(in[290] ^ in[632]); 
    assign layer_0[600] = in[978] & ~in[1009]; 
    assign layer_0[601] = in[316] & ~in[917]; 
    assign layer_0[602] = ~in[207]; 
    assign layer_0[603] = ~(in[483] ^ in[851]); 
    assign layer_0[604] = ~(in[596] & in[428]); 
    assign layer_0[605] = ~in[682] | (in[308] & in[682]); 
    assign layer_0[606] = ~in[872] | (in[872] & in[204]); 
    assign layer_0[607] = ~in[556] | (in[2] & in[556]); 
    assign layer_0[608] = in[173] & ~in[762]; 
    assign layer_0[609] = 1'b1; 
    assign layer_0[610] = in[46] ^ in[604]; 
    assign layer_0[611] = in[989] & in[554]; 
    assign layer_0[612] = in[1000] ^ in[999]; 
    assign layer_0[613] = in[478] ^ in[504]; 
    assign layer_0[614] = ~(in[477] ^ in[819]); 
    assign layer_0[615] = in[588] ^ in[483]; 
    assign layer_0[616] = ~(in[823] | in[599]); 
    assign layer_0[617] = ~(in[726] ^ in[384]); 
    assign layer_0[618] = in[841] & ~in[615]; 
    assign layer_0[619] = ~(in[384] ^ in[257]); 
    assign layer_0[620] = in[810] ^ in[701]; 
    assign layer_0[621] = ~in[180] | (in[180] & in[2]); 
    assign layer_0[622] = in[50] ^ in[852]; 
    assign layer_0[623] = ~(in[109] ^ in[210]); 
    assign layer_0[624] = in[533] | in[548]; 
    assign layer_0[625] = in[304] | in[1001]; 
    assign layer_0[626] = ~in[689]; 
    assign layer_0[627] = ~(in[491] & in[415]); 
    assign layer_0[628] = ~(in[56] ^ in[607]); 
    assign layer_0[629] = ~(in[538] | in[316]); 
    assign layer_0[630] = in[302] ^ in[713]; 
    assign layer_0[631] = in[719] & ~in[485]; 
    assign layer_0[632] = in[841] ^ in[940]; 
    assign layer_0[633] = in[885]; 
    assign layer_0[634] = in[84] & ~in[791]; 
    assign layer_0[635] = in[365] ^ in[837]; 
    assign layer_0[636] = in[104] & ~in[838]; 
    assign layer_0[637] = in[221] ^ in[488]; 
    assign layer_0[638] = in[920] ^ in[888]; 
    assign layer_0[639] = ~(in[333] | in[47]); 
    assign layer_0[640] = ~(in[253] ^ in[756]); 
    assign layer_0[641] = in[187] ^ in[873]; 
    assign layer_0[642] = ~(in[710] & in[635]); 
    assign layer_0[643] = ~in[546] | (in[72] & in[546]); 
    assign layer_0[644] = ~in[910]; 
    assign layer_0[645] = ~(in[484] & in[826]); 
    assign layer_0[646] = in[19] & ~in[868]; 
    assign layer_0[647] = ~(in[451] & in[8]); 
    assign layer_0[648] = ~(in[46] ^ in[744]); 
    assign layer_0[649] = in[66]; 
    assign layer_0[650] = in[600] ^ in[618]; 
    assign layer_0[651] = ~(in[465] ^ in[566]); 
    assign layer_0[652] = in[794] ^ in[823]; 
    assign layer_0[653] = 1'b1; 
    assign layer_0[654] = ~in[1016]; 
    assign layer_0[655] = ~in[312]; 
    assign layer_0[656] = in[594] ^ in[315]; 
    assign layer_0[657] = in[809] ^ in[639]; 
    assign layer_0[658] = in[401] ^ in[388]; 
    assign layer_0[659] = ~(in[119] & in[315]); 
    assign layer_0[660] = in[216] & in[984]; 
    assign layer_0[661] = in[425] | in[475]; 
    assign layer_0[662] = in[966] | in[436]; 
    assign layer_0[663] = ~(in[311] ^ in[264]); 
    assign layer_0[664] = in[30] | in[190]; 
    assign layer_0[665] = ~in[77] | (in[77] & in[808]); 
    assign layer_0[666] = in[704] ^ in[307]; 
    assign layer_0[667] = in[267] | in[338]; 
    assign layer_0[668] = ~(in[852] ^ in[936]); 
    assign layer_0[669] = ~(in[786] | in[888]); 
    assign layer_0[670] = ~in[146] | (in[930] & in[146]); 
    assign layer_0[671] = ~in[101] | (in[494] & in[101]); 
    assign layer_0[672] = ~(in[628] ^ in[189]); 
    assign layer_0[673] = in[517] ^ in[838]; 
    assign layer_0[674] = in[954] ^ in[467]; 
    assign layer_0[675] = ~(in[884] ^ in[996]); 
    assign layer_0[676] = ~(in[518] | in[667]); 
    assign layer_0[677] = ~in[566]; 
    assign layer_0[678] = in[205]; 
    assign layer_0[679] = ~(in[868] ^ in[261]); 
    assign layer_0[680] = ~(in[833] | in[352]); 
    assign layer_0[681] = in[459] | in[817]; 
    assign layer_0[682] = in[865] ^ in[583]; 
    assign layer_0[683] = ~(in[264] ^ in[266]); 
    assign layer_0[684] = ~(in[617] & in[679]); 
    assign layer_0[685] = ~(in[411] ^ in[790]); 
    assign layer_0[686] = in[277]; 
    assign layer_0[687] = ~(in[347] & in[356]); 
    assign layer_0[688] = ~in[519] | (in[982] & in[519]); 
    assign layer_0[689] = ~(in[945] | in[77]); 
    assign layer_0[690] = in[809] ^ in[677]; 
    assign layer_0[691] = ~in[600] | (in[600] & in[834]); 
    assign layer_0[692] = ~(in[505] ^ in[507]); 
    assign layer_0[693] = in[311] & in[35]; 
    assign layer_0[694] = in[413] ^ in[741]; 
    assign layer_0[695] = ~in[954] | (in[565] & in[954]); 
    assign layer_0[696] = ~in[82]; 
    assign layer_0[697] = in[892] & ~in[741]; 
    assign layer_0[698] = ~in[803] | (in[803] & in[722]); 
    assign layer_0[699] = ~in[433]; 
    assign layer_0[700] = ~in[614] | (in[614] & in[465]); 
    assign layer_0[701] = in[886] ^ in[926]; 
    assign layer_0[702] = in[55] ^ in[904]; 
    assign layer_0[703] = in[930] ^ in[357]; 
    assign layer_0[704] = in[253] ^ in[746]; 
    assign layer_0[705] = ~(in[776] ^ in[83]); 
    assign layer_0[706] = ~in[1013] | (in[1013] & in[931]); 
    assign layer_0[707] = in[939] ^ in[937]; 
    assign layer_0[708] = ~in[98] | (in[98] & in[221]); 
    assign layer_0[709] = in[874] ^ in[90]; 
    assign layer_0[710] = ~(in[191] ^ in[944]); 
    assign layer_0[711] = ~(in[280] ^ in[549]); 
    assign layer_0[712] = ~in[603]; 
    assign layer_0[713] = in[160]; 
    assign layer_0[714] = in[635]; 
    assign layer_0[715] = ~(in[204] & in[72]); 
    assign layer_0[716] = in[221] | in[853]; 
    assign layer_0[717] = in[146]; 
    assign layer_0[718] = ~in[96] | (in[57] & in[96]); 
    assign layer_0[719] = ~(in[69] | in[535]); 
    assign layer_0[720] = ~(in[807] ^ in[299]); 
    assign layer_0[721] = ~in[252] | (in[777] & in[252]); 
    assign layer_0[722] = ~in[664] | (in[290] & in[664]); 
    assign layer_0[723] = in[905] & ~in[550]; 
    assign layer_0[724] = in[822] ^ in[684]; 
    assign layer_0[725] = in[553] & in[584]; 
    assign layer_0[726] = ~(in[441] ^ in[30]); 
    assign layer_0[727] = in[54] & in[82]; 
    assign layer_0[728] = in[843]; 
    assign layer_0[729] = ~(in[353] ^ in[824]); 
    assign layer_0[730] = ~in[473] | (in[535] & in[473]); 
    assign layer_0[731] = 1'b0; 
    assign layer_0[732] = in[317] ^ in[587]; 
    assign layer_0[733] = ~in[868]; 
    assign layer_0[734] = ~(in[668] | in[1017]); 
    assign layer_0[735] = ~(in[591] & in[359]); 
    assign layer_0[736] = ~in[300] | (in[300] & in[794]); 
    assign layer_0[737] = in[667]; 
    assign layer_0[738] = ~in[617] | (in[617] & in[252]); 
    assign layer_0[739] = in[486] & ~in[784]; 
    assign layer_0[740] = in[204] & ~in[387]; 
    assign layer_0[741] = in[939] ^ in[908]; 
    assign layer_0[742] = in[93] ^ in[935]; 
    assign layer_0[743] = 1'b1; 
    assign layer_0[744] = ~in[948] | (in[958] & in[948]); 
    assign layer_0[745] = in[724]; 
    assign layer_0[746] = ~in[72]; 
    assign layer_0[747] = ~(in[990] | in[374]); 
    assign layer_0[748] = in[264]; 
    assign layer_0[749] = ~(in[465] & in[55]); 
    assign layer_0[750] = in[643]; 
    assign layer_0[751] = in[241] & ~in[283]; 
    assign layer_0[752] = ~(in[631] ^ in[940]); 
    assign layer_0[753] = in[243] & ~in[446]; 
    assign layer_0[754] = in[436] ^ in[252]; 
    assign layer_0[755] = in[596] ^ in[857]; 
    assign layer_0[756] = ~in[986] | (in[968] & in[986]); 
    assign layer_0[757] = in[1004] & ~in[758]; 
    assign layer_0[758] = in[29] ^ in[129]; 
    assign layer_0[759] = ~in[422] | (in[422] & in[850]); 
    assign layer_0[760] = ~in[837]; 
    assign layer_0[761] = ~in[844]; 
    assign layer_0[762] = in[607]; 
    assign layer_0[763] = ~(in[162] | in[177]); 
    assign layer_0[764] = in[868]; 
    assign layer_0[765] = ~(in[4] ^ in[826]); 
    assign layer_0[766] = in[457]; 
    assign layer_0[767] = ~in[931] | (in[931] & in[657]); 
    assign layer_0[768] = ~(in[241] ^ in[987]); 
    assign layer_0[769] = ~in[215] | (in[573] & in[215]); 
    assign layer_0[770] = ~(in[414] & in[856]); 
    assign layer_0[771] = ~(in[477] ^ in[14]); 
    assign layer_0[772] = in[838] ^ in[837]; 
    assign layer_0[773] = ~in[118] | (in[629] & in[118]); 
    assign layer_0[774] = in[265] & ~in[588]; 
    assign layer_0[775] = 1'b1; 
    assign layer_0[776] = ~in[282] | (in[282] & in[967]); 
    assign layer_0[777] = in[636] ^ in[702]; 
    assign layer_0[778] = in[938] ^ in[317]; 
    assign layer_0[779] = ~in[373] | (in[373] & in[254]); 
    assign layer_0[780] = in[634] & ~in[568]; 
    assign layer_0[781] = in[99] ^ in[842]; 
    assign layer_0[782] = in[286] | in[342]; 
    assign layer_0[783] = ~(in[738] | in[901]); 
    assign layer_0[784] = in[498]; 
    assign layer_0[785] = in[371]; 
    assign layer_0[786] = in[565] | in[598]; 
    assign layer_0[787] = ~(in[265] ^ in[96]); 
    assign layer_0[788] = in[605] & in[99]; 
    assign layer_0[789] = ~(in[629] & in[743]); 
    assign layer_0[790] = ~in[8] | (in[8] & in[1015]); 
    assign layer_0[791] = in[339] ^ in[460]; 
    assign layer_0[792] = in[603] & in[660]; 
    assign layer_0[793] = in[122] & ~in[955]; 
    assign layer_0[794] = ~(in[695] | in[432]); 
    assign layer_0[795] = in[35] ^ in[845]; 
    assign layer_0[796] = ~(in[525] & in[466]); 
    assign layer_0[797] = ~(in[838] ^ in[842]); 
    assign layer_0[798] = in[411] & in[467]; 
    assign layer_0[799] = ~(in[690] & in[949]); 
    assign layer_0[800] = in[917] & ~in[596]; 
    assign layer_0[801] = ~in[234] | (in[807] & in[234]); 
    assign layer_0[802] = in[839] | in[868]; 
    assign layer_0[803] = in[278]; 
    assign layer_0[804] = ~(in[855] ^ in[348]); 
    assign layer_0[805] = ~(in[564] ^ in[19]); 
    assign layer_0[806] = ~(in[931] ^ in[808]); 
    assign layer_0[807] = ~(in[596] | in[880]); 
    assign layer_0[808] = in[681]; 
    assign layer_0[809] = in[557] | in[764]; 
    assign layer_0[810] = in[997] ^ in[142]; 
    assign layer_0[811] = ~(in[509] & in[204]); 
    assign layer_0[812] = ~(in[795] ^ in[651]); 
    assign layer_0[813] = ~(in[488] & in[227]); 
    assign layer_0[814] = 1'b0; 
    assign layer_0[815] = in[614] & ~in[354]; 
    assign layer_0[816] = ~in[899]; 
    assign layer_0[817] = ~in[874]; 
    assign layer_0[818] = in[957] & ~in[916]; 
    assign layer_0[819] = ~in[757]; 
    assign layer_0[820] = in[861] ^ in[294]; 
    assign layer_0[821] = ~in[411]; 
    assign layer_0[822] = 1'b0; 
    assign layer_0[823] = ~(in[897] | in[185]); 
    assign layer_0[824] = ~(in[602] & in[244]); 
    assign layer_0[825] = in[33]; 
    assign layer_0[826] = ~(in[161] ^ in[808]); 
    assign layer_0[827] = in[7]; 
    assign layer_0[828] = in[368]; 
    assign layer_0[829] = in[765]; 
    assign layer_0[830] = in[956] ^ in[487]; 
    assign layer_0[831] = ~in[459] | (in[548] & in[459]); 
    assign layer_0[832] = in[279]; 
    assign layer_0[833] = ~(in[99] ^ in[226]); 
    assign layer_0[834] = in[614] ^ in[266]; 
    assign layer_0[835] = ~(in[78] ^ in[276]); 
    assign layer_0[836] = ~in[412] | (in[412] & in[96]); 
    assign layer_0[837] = in[946] & ~in[114]; 
    assign layer_0[838] = in[600] & ~in[871]; 
    assign layer_0[839] = in[932] | in[855]; 
    assign layer_0[840] = ~in[485] | (in[485] & in[943]); 
    assign layer_0[841] = ~in[727]; 
    assign layer_0[842] = in[537] & ~in[462]; 
    assign layer_0[843] = in[625]; 
    assign layer_0[844] = in[255] & ~in[904]; 
    assign layer_0[845] = ~in[71] | (in[71] & in[67]); 
    assign layer_0[846] = ~(in[341] | in[489]); 
    assign layer_0[847] = ~(in[374] | in[837]); 
    assign layer_0[848] = ~(in[84] ^ in[447]); 
    assign layer_0[849] = in[845] & in[116]; 
    assign layer_0[850] = ~in[972]; 
    assign layer_0[851] = in[360] & ~in[746]; 
    assign layer_0[852] = in[622] ^ in[603]; 
    assign layer_0[853] = ~(in[692] | in[660]); 
    assign layer_0[854] = in[602] & ~in[1011]; 
    assign layer_0[855] = ~in[876]; 
    assign layer_0[856] = in[994] & in[710]; 
    assign layer_0[857] = ~(in[877] & in[388]); 
    assign layer_0[858] = ~(in[627] ^ in[907]); 
    assign layer_0[859] = in[174]; 
    assign layer_0[860] = in[952] & ~in[509]; 
    assign layer_0[861] = in[261] & ~in[725]; 
    assign layer_0[862] = ~(in[568] ^ in[569]); 
    assign layer_0[863] = ~(in[938] ^ in[67]); 
    assign layer_0[864] = ~in[874]; 
    assign layer_0[865] = ~in[773] | (in[683] & in[773]); 
    assign layer_0[866] = ~in[308]; 
    assign layer_0[867] = ~(in[1000] ^ in[808]); 
    assign layer_0[868] = in[419] & ~in[839]; 
    assign layer_0[869] = ~in[842] | (in[429] & in[842]); 
    assign layer_0[870] = in[468] | in[955]; 
    assign layer_0[871] = ~(in[892] ^ in[943]); 
    assign layer_0[872] = in[430] ^ in[809]; 
    assign layer_0[873] = ~in[651]; 
    assign layer_0[874] = ~in[2]; 
    assign layer_0[875] = ~in[191] | (in[191] & in[68]); 
    assign layer_0[876] = 1'b0; 
    assign layer_0[877] = in[63] ^ in[189]; 
    assign layer_0[878] = in[466] ^ in[569]; 
    assign layer_0[879] = ~in[505]; 
    assign layer_0[880] = ~in[568] | (in[295] & in[568]); 
    assign layer_0[881] = ~(in[201] ^ in[871]); 
    assign layer_0[882] = in[171] & in[377]; 
    assign layer_0[883] = ~in[176]; 
    assign layer_0[884] = ~in[793]; 
    assign layer_0[885] = ~(in[5] & in[920]); 
    assign layer_0[886] = in[580] & ~in[349]; 
    assign layer_0[887] = ~(in[156] ^ in[919]); 
    assign layer_0[888] = ~in[8] | (in[856] & in[8]); 
    assign layer_0[889] = ~in[368] | (in[368] & in[498]); 
    assign layer_0[890] = ~(in[493] | in[674]); 
    assign layer_0[891] = ~(in[987] ^ in[588]); 
    assign layer_0[892] = in[951] ^ in[875]; 
    assign layer_0[893] = in[595] & ~in[776]; 
    assign layer_0[894] = ~(in[775] | in[618]); 
    assign layer_0[895] = ~(in[692] ^ in[227]); 
    assign layer_0[896] = in[931] & ~in[78]; 
    assign layer_0[897] = ~(in[447] ^ in[84]); 
    assign layer_0[898] = in[549] | in[555]; 
    assign layer_0[899] = in[302] ^ in[450]; 
    assign layer_0[900] = in[264] | in[494]; 
    assign layer_0[901] = in[267] | in[111]; 
    assign layer_0[902] = in[322] ^ in[77]; 
    assign layer_0[903] = in[267] | in[274]; 
    assign layer_0[904] = in[953] ^ in[42]; 
    assign layer_0[905] = ~(in[804] ^ in[924]); 
    assign layer_0[906] = ~(in[674] & in[291]); 
    assign layer_0[907] = ~(in[871] ^ in[912]); 
    assign layer_0[908] = in[131] | in[673]; 
    assign layer_0[909] = in[940] ^ in[59]; 
    assign layer_0[910] = ~(in[515] ^ in[1016]); 
    assign layer_0[911] = ~in[273]; 
    assign layer_0[912] = ~in[468] | (in[987] & in[468]); 
    assign layer_0[913] = ~in[972]; 
    assign layer_0[914] = in[246] & ~in[549]; 
    assign layer_0[915] = in[618] ^ in[603]; 
    assign layer_0[916] = in[989] ^ in[307]; 
    assign layer_0[917] = in[94] ^ in[462]; 
    assign layer_0[918] = ~in[161]; 
    assign layer_0[919] = in[660] & in[570]; 
    assign layer_0[920] = in[466] & in[621]; 
    assign layer_0[921] = ~(in[474] | in[338]); 
    assign layer_0[922] = ~(in[582] ^ in[807]); 
    assign layer_0[923] = in[227] & in[296]; 
    assign layer_0[924] = ~(in[276] ^ in[115]); 
    assign layer_0[925] = in[76] & ~in[600]; 
    assign layer_0[926] = in[871] & ~in[44]; 
    assign layer_0[927] = in[87]; 
    assign layer_0[928] = in[1017]; 
    assign layer_0[929] = in[176] & in[662]; 
    assign layer_0[930] = in[933] ^ in[249]; 
    assign layer_0[931] = in[297] & ~in[17]; 
    assign layer_0[932] = in[934] & ~in[29]; 
    assign layer_0[933] = ~(in[917] ^ in[934]); 
    assign layer_0[934] = ~(in[46] | in[421]); 
    assign layer_0[935] = ~(in[596] ^ in[843]); 
    assign layer_0[936] = ~(in[508] | in[18]); 
    assign layer_0[937] = in[975]; 
    assign layer_0[938] = ~(in[971] ^ in[747]); 
    assign layer_0[939] = in[876] ^ in[96]; 
    assign layer_0[940] = in[649] & ~in[451]; 
    assign layer_0[941] = ~(in[203] ^ in[610]); 
    assign layer_0[942] = in[2] & in[105]; 
    assign layer_0[943] = in[476] ^ in[762]; 
    assign layer_0[944] = in[317] ^ in[533]; 
    assign layer_0[945] = in[682] & ~in[766]; 
    assign layer_0[946] = ~in[183] | (in[563] & in[183]); 
    assign layer_0[947] = ~(in[730] ^ in[658]); 
    assign layer_0[948] = in[413] & ~in[492]; 
    assign layer_0[949] = in[688] & in[473]; 
    assign layer_0[950] = ~in[939] | (in[980] & in[939]); 
    assign layer_0[951] = ~(in[238] ^ in[687]); 
    assign layer_0[952] = in[922] ^ in[85]; 
    assign layer_0[953] = in[936] ^ in[937]; 
    assign layer_0[954] = ~(in[588] ^ in[581]); 
    assign layer_0[955] = in[419] | in[1022]; 
    assign layer_0[956] = ~in[436] | (in[436] & in[732]); 
    assign layer_0[957] = ~in[131] | (in[467] & in[131]); 
    assign layer_0[958] = in[306]; 
    assign layer_0[959] = 1'b0; 
    assign layer_0[960] = ~in[859] | (in[859] & in[598]); 
    assign layer_0[961] = in[1001] ^ in[627]; 
    assign layer_0[962] = 1'b1; 
    assign layer_0[963] = ~in[439] | (in[439] & in[822]); 
    assign layer_0[964] = in[708] ^ in[757]; 
    assign layer_0[965] = ~(in[319] ^ in[296]); 
    assign layer_0[966] = in[732] ^ in[907]; 
    assign layer_0[967] = ~(in[3] | in[606]); 
    assign layer_0[968] = in[82] ^ in[673]; 
    assign layer_0[969] = ~in[982] | (in[982] & in[708]); 
    assign layer_0[970] = ~(in[865] | in[873]); 
    assign layer_0[971] = ~(in[53] & in[852]); 
    assign layer_0[972] = in[281] ^ in[252]; 
    assign layer_0[973] = ~(in[995] | in[275]); 
    assign layer_0[974] = ~in[26] | (in[800] & in[26]); 
    assign layer_0[975] = in[776] ^ in[83]; 
    assign layer_0[976] = ~in[243]; 
    assign layer_0[977] = ~in[844] | (in[578] & in[844]); 
    assign layer_0[978] = ~in[230] | (in[554] & in[230]); 
    assign layer_0[979] = in[967] ^ in[570]; 
    assign layer_0[980] = in[533] ^ in[44]; 
    assign layer_0[981] = ~in[905] | (in[808] & in[905]); 
    assign layer_0[982] = ~in[371]; 
    assign layer_0[983] = in[775] ^ in[532]; 
    assign layer_0[984] = in[883] | in[253]; 
    assign layer_0[985] = in[808] ^ in[473]; 
    assign layer_0[986] = ~(in[607] ^ in[844]); 
    assign layer_0[987] = in[151] ^ in[126]; 
    assign layer_0[988] = in[499] | in[363]; 
    assign layer_0[989] = in[987] ^ in[776]; 
    assign layer_0[990] = in[253] & in[37]; 
    assign layer_0[991] = in[809] ^ in[351]; 
    assign layer_0[992] = in[496] | in[278]; 
    assign layer_0[993] = ~in[164] | (in[164] & in[1001]); 
    assign layer_0[994] = in[427]; 
    assign layer_0[995] = ~(in[562] ^ in[794]); 
    assign layer_0[996] = in[774] & ~in[984]; 
    assign layer_0[997] = ~(in[62] | in[248]); 
    assign layer_0[998] = in[1017] ^ in[612]; 
    assign layer_0[999] = ~(in[933] ^ in[713]); 
    assign layer_0[1000] = ~in[857] | (in[178] & in[857]); 
    assign layer_0[1001] = ~in[143] | (in[143] & in[948]); 
    assign layer_0[1002] = ~(in[302] ^ in[905]); 
    assign layer_0[1003] = ~(in[875] ^ in[982]); 
    assign layer_0[1004] = in[590] & in[73]; 
    assign layer_0[1005] = ~(in[345] | in[547]); 
    assign layer_0[1006] = in[461] ^ in[316]; 
    assign layer_0[1007] = in[291]; 
    assign layer_0[1008] = in[276] ^ in[434]; 
    assign layer_0[1009] = in[918] ^ in[870]; 
    assign layer_0[1010] = in[893] ^ in[62]; 
    assign layer_0[1011] = ~in[1015]; 
    assign layer_0[1012] = in[660] ^ in[859]; 
    assign layer_0[1013] = in[906] | in[422]; 
    assign layer_0[1014] = in[865] & in[104]; 
    assign layer_0[1015] = ~in[437] | (in[437] & in[20]); 
    assign layer_0[1016] = ~in[128] | (in[128] & in[62]); 
    assign layer_0[1017] = ~in[375] | (in[375] & in[875]); 
    assign layer_0[1018] = in[724] ^ in[454]; 
    assign layer_0[1019] = in[60] ^ in[42]; 
    assign layer_0[1020] = ~(in[1016] | in[686]); 
    assign layer_0[1021] = ~in[29]; 
    assign layer_0[1022] = ~(in[435] ^ in[684]); 
    assign layer_0[1023] = ~in[50]; 
    assign layer_0[1024] = in[905] & in[549]; 
    assign layer_0[1025] = in[835] ^ in[802]; 
    assign layer_0[1026] = ~in[342] | (in[488] & in[342]); 
    assign layer_0[1027] = ~(in[356] & in[413]); 
    assign layer_0[1028] = ~in[445] | (in[445] & in[310]); 
    assign layer_0[1029] = ~in[743] | (in[826] & in[743]); 
    assign layer_0[1030] = in[931] & in[765]; 
    assign layer_0[1031] = in[110]; 
    assign layer_0[1032] = in[436]; 
    assign layer_0[1033] = in[989] ^ in[654]; 
    assign layer_0[1034] = in[621] & in[694]; 
    assign layer_0[1035] = in[948] & ~in[794]; 
    assign layer_0[1036] = ~(in[902] ^ in[126]); 
    assign layer_0[1037] = ~(in[323] ^ in[460]); 
    assign layer_0[1038] = in[69] & ~in[536]; 
    assign layer_0[1039] = in[600]; 
    assign layer_0[1040] = in[1013] | in[821]; 
    assign layer_0[1041] = ~in[52] | (in[379] & in[52]); 
    assign layer_0[1042] = ~in[984]; 
    assign layer_0[1043] = ~(in[952] ^ in[76]); 
    assign layer_0[1044] = ~(in[973] | in[96]); 
    assign layer_0[1045] = in[225] & ~in[989]; 
    assign layer_0[1046] = ~(in[811] & in[222]); 
    assign layer_0[1047] = ~in[325]; 
    assign layer_0[1048] = in[417] & ~in[593]; 
    assign layer_0[1049] = in[608] | in[471]; 
    assign layer_0[1050] = ~in[685]; 
    assign layer_0[1051] = in[824] | in[828]; 
    assign layer_0[1052] = ~in[857] | (in[857] & in[859]); 
    assign layer_0[1053] = ~in[647] | (in[352] & in[647]); 
    assign layer_0[1054] = ~(in[276] ^ in[291]); 
    assign layer_0[1055] = in[997] | in[855]; 
    assign layer_0[1056] = in[22] & ~in[843]; 
    assign layer_0[1057] = in[986] ^ in[920]; 
    assign layer_0[1058] = ~(in[827] ^ in[714]); 
    assign layer_0[1059] = ~(in[406] ^ in[884]); 
    assign layer_0[1060] = ~(in[716] ^ in[844]); 
    assign layer_0[1061] = in[1016] | in[412]; 
    assign layer_0[1062] = in[869] ^ in[537]; 
    assign layer_0[1063] = in[474] & ~in[234]; 
    assign layer_0[1064] = in[462] ^ in[193]; 
    assign layer_0[1065] = ~(in[171] ^ in[281]); 
    assign layer_0[1066] = ~(in[873] ^ in[264]); 
    assign layer_0[1067] = ~in[731] | (in[731] & in[451]); 
    assign layer_0[1068] = ~(in[636] & in[60]); 
    assign layer_0[1069] = ~in[548]; 
    assign layer_0[1070] = ~(in[1020] | in[622]); 
    assign layer_0[1071] = in[579] ^ in[612]; 
    assign layer_0[1072] = ~in[325]; 
    assign layer_0[1073] = ~in[708] | (in[340] & in[708]); 
    assign layer_0[1074] = in[749] ^ in[907]; 
    assign layer_0[1075] = ~(in[477] & in[466]); 
    assign layer_0[1076] = ~in[899]; 
    assign layer_0[1077] = ~(in[451] ^ in[983]); 
    assign layer_0[1078] = in[597] & ~in[270]; 
    assign layer_0[1079] = in[730] & in[536]; 
    assign layer_0[1080] = in[712] & in[410]; 
    assign layer_0[1081] = ~(in[353] ^ in[804]); 
    assign layer_0[1082] = ~(in[111] ^ in[445]); 
    assign layer_0[1083] = in[502] | in[714]; 
    assign layer_0[1084] = ~(in[50] & in[551]); 
    assign layer_0[1085] = ~(in[262] ^ in[238]); 
    assign layer_0[1086] = ~in[268]; 
    assign layer_0[1087] = in[508]; 
    assign layer_0[1088] = ~(in[903] ^ in[114]); 
    assign layer_0[1089] = ~in[434] | (in[434] & in[954]); 
    assign layer_0[1090] = ~in[316]; 
    assign layer_0[1091] = 1'b1; 
    assign layer_0[1092] = ~in[67] | (in[67] & in[80]); 
    assign layer_0[1093] = ~(in[232] & in[620]); 
    assign layer_0[1094] = in[705] ^ in[22]; 
    assign layer_0[1095] = in[910] ^ in[952]; 
    assign layer_0[1096] = ~(in[470] ^ in[125]); 
    assign layer_0[1097] = ~(in[567] ^ in[307]); 
    assign layer_0[1098] = in[268] ^ in[301]; 
    assign layer_0[1099] = in[53] ^ in[915]; 
    assign layer_0[1100] = ~(in[616] ^ in[667]); 
    assign layer_0[1101] = ~(in[319] ^ in[914]); 
    assign layer_0[1102] = in[581]; 
    assign layer_0[1103] = in[427] ^ in[707]; 
    assign layer_0[1104] = in[894] & ~in[299]; 
    assign layer_0[1105] = in[761] ^ in[968]; 
    assign layer_0[1106] = ~in[559] | (in[82] & in[559]); 
    assign layer_0[1107] = ~in[99]; 
    assign layer_0[1108] = ~(in[1015] ^ in[1016]); 
    assign layer_0[1109] = in[271]; 
    assign layer_0[1110] = ~(in[276] ^ in[981]); 
    assign layer_0[1111] = ~in[129]; 
    assign layer_0[1112] = ~(in[50] ^ in[483]); 
    assign layer_0[1113] = ~(in[648] ^ in[649]); 
    assign layer_0[1114] = ~in[98] | (in[808] & in[98]); 
    assign layer_0[1115] = ~in[920] | (in[115] & in[920]); 
    assign layer_0[1116] = ~in[552] | (in[775] & in[552]); 
    assign layer_0[1117] = ~(in[824] ^ in[507]); 
    assign layer_0[1118] = ~(in[903] ^ in[901]); 
    assign layer_0[1119] = in[595] & ~in[998]; 
    assign layer_0[1120] = ~(in[392] ^ in[284]); 
    assign layer_0[1121] = in[913] ^ in[100]; 
    assign layer_0[1122] = ~(in[552] & in[899]); 
    assign layer_0[1123] = in[645] ^ in[630]; 
    assign layer_0[1124] = ~(in[859] ^ in[518]); 
    assign layer_0[1125] = in[269] & ~in[336]; 
    assign layer_0[1126] = in[661]; 
    assign layer_0[1127] = in[236] & in[56]; 
    assign layer_0[1128] = in[295] & ~in[30]; 
    assign layer_0[1129] = in[879]; 
    assign layer_0[1130] = ~(in[647] ^ in[918]); 
    assign layer_0[1131] = ~in[928]; 
    assign layer_0[1132] = ~(in[509] ^ in[997]); 
    assign layer_0[1133] = ~(in[552] ^ in[98]); 
    assign layer_0[1134] = in[299] & ~in[741]; 
    assign layer_0[1135] = ~(in[547] ^ in[611]); 
    assign layer_0[1136] = ~(in[820] | in[895]); 
    assign layer_0[1137] = in[790] ^ in[690]; 
    assign layer_0[1138] = in[61] & ~in[795]; 
    assign layer_0[1139] = in[966] & ~in[554]; 
    assign layer_0[1140] = ~(in[102] ^ in[940]); 
    assign layer_0[1141] = ~(in[723] ^ in[170]); 
    assign layer_0[1142] = in[922]; 
    assign layer_0[1143] = ~in[646] | (in[572] & in[646]); 
    assign layer_0[1144] = ~in[872]; 
    assign layer_0[1145] = in[215] | in[196]; 
    assign layer_0[1146] = ~in[953]; 
    assign layer_0[1147] = ~(in[686] ^ in[882]); 
    assign layer_0[1148] = in[554]; 
    assign layer_0[1149] = in[49] ^ in[383]; 
    assign layer_0[1150] = in[649] & in[714]; 
    assign layer_0[1151] = ~(in[122] ^ in[200]); 
    assign layer_0[1152] = in[734] ^ in[729]; 
    assign layer_0[1153] = ~(in[929] | in[254]); 
    assign layer_0[1154] = ~in[333] | (in[182] & in[333]); 
    assign layer_0[1155] = ~(in[643] ^ in[668]); 
    assign layer_0[1156] = in[383] | in[818]; 
    assign layer_0[1157] = ~in[723]; 
    assign layer_0[1158] = in[261] ^ in[825]; 
    assign layer_0[1159] = in[588] & ~in[476]; 
    assign layer_0[1160] = ~(in[858] ^ in[873]); 
    assign layer_0[1161] = ~(in[43] ^ in[56]); 
    assign layer_0[1162] = in[844] ^ in[46]; 
    assign layer_0[1163] = in[571] & ~in[268]; 
    assign layer_0[1164] = in[635] & ~in[658]; 
    assign layer_0[1165] = in[892]; 
    assign layer_0[1166] = ~in[156] | (in[156] & in[573]); 
    assign layer_0[1167] = in[920] ^ in[808]; 
    assign layer_0[1168] = in[903]; 
    assign layer_0[1169] = in[52]; 
    assign layer_0[1170] = ~in[872] | (in[547] & in[872]); 
    assign layer_0[1171] = ~in[611] | (in[865] & in[611]); 
    assign layer_0[1172] = in[55] & ~in[320]; 
    assign layer_0[1173] = ~(in[263] ^ in[356]); 
    assign layer_0[1174] = ~(in[93] ^ in[875]); 
    assign layer_0[1175] = ~in[907] | (in[843] & in[907]); 
    assign layer_0[1176] = in[588] | in[914]; 
    assign layer_0[1177] = in[572] & in[300]; 
    assign layer_0[1178] = in[851] ^ in[64]; 
    assign layer_0[1179] = ~in[871] | (in[871] & in[93]); 
    assign layer_0[1180] = in[664] & in[978]; 
    assign layer_0[1181] = in[195] ^ in[793]; 
    assign layer_0[1182] = in[373] & in[25]; 
    assign layer_0[1183] = ~(in[984] ^ in[794]); 
    assign layer_0[1184] = ~(in[18] | in[317]); 
    assign layer_0[1185] = ~(in[604] ^ in[568]); 
    assign layer_0[1186] = ~(in[849] & in[380]); 
    assign layer_0[1187] = ~in[913] | (in[913] & in[178]); 
    assign layer_0[1188] = ~in[852]; 
    assign layer_0[1189] = in[276] ^ in[146]; 
    assign layer_0[1190] = ~(in[687] ^ in[342]); 
    assign layer_0[1191] = in[636]; 
    assign layer_0[1192] = ~(in[269] ^ in[572]); 
    assign layer_0[1193] = ~in[966] | (in[49] & in[966]); 
    assign layer_0[1194] = in[294] & ~in[376]; 
    assign layer_0[1195] = in[661] ^ in[162]; 
    assign layer_0[1196] = 1'b0; 
    assign layer_0[1197] = in[875] | in[622]; 
    assign layer_0[1198] = in[460] ^ in[895]; 
    assign layer_0[1199] = in[929] & ~in[953]; 
    assign layer_0[1200] = ~in[603] | (in[603] & in[225]); 
    assign layer_0[1201] = in[224] & ~in[82]; 
    assign layer_0[1202] = in[352]; 
    assign layer_0[1203] = ~(in[206] ^ in[366]); 
    assign layer_0[1204] = 1'b0; 
    assign layer_0[1205] = in[983] & ~in[623]; 
    assign layer_0[1206] = ~in[546] | (in[546] & in[436]); 
    assign layer_0[1207] = ~in[262]; 
    assign layer_0[1208] = ~(in[949] ^ in[98]); 
    assign layer_0[1209] = ~in[504]; 
    assign layer_0[1210] = ~in[648]; 
    assign layer_0[1211] = ~in[81]; 
    assign layer_0[1212] = ~in[53] | (in[53] & in[544]); 
    assign layer_0[1213] = in[325] ^ in[897]; 
    assign layer_0[1214] = ~in[146] | (in[944] & in[146]); 
    assign layer_0[1215] = 1'b1; 
    assign layer_0[1216] = ~(in[950] ^ in[871]); 
    assign layer_0[1217] = ~(in[700] ^ in[989]); 
    assign layer_0[1218] = ~in[587] | (in[587] & in[265]); 
    assign layer_0[1219] = in[968] & in[617]; 
    assign layer_0[1220] = in[169] & ~in[1002]; 
    assign layer_0[1221] = in[972] ^ in[86]; 
    assign layer_0[1222] = in[280]; 
    assign layer_0[1223] = in[837] ^ in[66]; 
    assign layer_0[1224] = ~(in[850] ^ in[537]); 
    assign layer_0[1225] = ~(in[775] ^ in[244]); 
    assign layer_0[1226] = ~(in[267] ^ in[508]); 
    assign layer_0[1227] = ~(in[997] ^ in[990]); 
    assign layer_0[1228] = in[51]; 
    assign layer_0[1229] = in[644] & in[314]; 
    assign layer_0[1230] = in[689]; 
    assign layer_0[1231] = in[58] ^ in[951]; 
    assign layer_0[1232] = ~(in[792] ^ in[12]); 
    assign layer_0[1233] = in[858]; 
    assign layer_0[1234] = ~in[953]; 
    assign layer_0[1235] = in[613]; 
    assign layer_0[1236] = ~(in[202] & in[691]); 
    assign layer_0[1237] = ~(in[12] ^ in[550]); 
    assign layer_0[1238] = ~(in[251] & in[986]); 
    assign layer_0[1239] = in[680] ^ in[698]; 
    assign layer_0[1240] = ~in[100]; 
    assign layer_0[1241] = ~(in[293] ^ in[971]); 
    assign layer_0[1242] = in[152] & ~in[98]; 
    assign layer_0[1243] = in[362] ^ in[67]; 
    assign layer_0[1244] = in[885] | in[60]; 
    assign layer_0[1245] = in[222] & ~in[276]; 
    assign layer_0[1246] = in[48] | in[477]; 
    assign layer_0[1247] = ~in[492] | (in[65] & in[492]); 
    assign layer_0[1248] = in[218] & in[571]; 
    assign layer_0[1249] = ~in[158] | (in[470] & in[158]); 
    assign layer_0[1250] = ~(in[862] ^ in[223]); 
    assign layer_0[1251] = in[576] & in[522]; 
    assign layer_0[1252] = ~(in[668] & in[402]); 
    assign layer_0[1253] = in[951]; 
    assign layer_0[1254] = ~(in[628] ^ in[924]); 
    assign layer_0[1255] = in[28] | in[370]; 
    assign layer_0[1256] = ~(in[12] ^ in[201]); 
    assign layer_0[1257] = in[995] | in[581]; 
    assign layer_0[1258] = ~(in[284] | in[588]); 
    assign layer_0[1259] = 1'b0; 
    assign layer_0[1260] = ~(in[318] | in[876]); 
    assign layer_0[1261] = ~in[412] | (in[412] & in[700]); 
    assign layer_0[1262] = in[504] ^ in[467]; 
    assign layer_0[1263] = ~(in[462] ^ in[804]); 
    assign layer_0[1264] = in[717] & ~in[988]; 
    assign layer_0[1265] = 1'b1; 
    assign layer_0[1266] = in[442] & ~in[74]; 
    assign layer_0[1267] = ~(in[628] ^ in[635]); 
    assign layer_0[1268] = ~(in[934] ^ in[951]); 
    assign layer_0[1269] = in[792] | in[809]; 
    assign layer_0[1270] = ~in[687] | (in[687] & in[643]); 
    assign layer_0[1271] = in[195] ^ in[456]; 
    assign layer_0[1272] = ~(in[913] | in[456]); 
    assign layer_0[1273] = in[365] & ~in[990]; 
    assign layer_0[1274] = ~(in[249] | in[958]); 
    assign layer_0[1275] = in[269] & in[859]; 
    assign layer_0[1276] = ~in[918] | (in[918] & in[876]); 
    assign layer_0[1277] = in[65] | in[898]; 
    assign layer_0[1278] = in[216] ^ in[1]; 
    assign layer_0[1279] = in[607]; 
    assign layer_0[1280] = in[509]; 
    assign layer_0[1281] = ~(in[888] ^ in[841]); 
    assign layer_0[1282] = ~in[402] | (in[435] & in[402]); 
    assign layer_0[1283] = in[34] & ~in[349]; 
    assign layer_0[1284] = ~(in[491] ^ in[728]); 
    assign layer_0[1285] = in[809] | in[567]; 
    assign layer_0[1286] = ~in[417] | (in[688] & in[417]); 
    assign layer_0[1287] = in[631] & ~in[890]; 
    assign layer_0[1288] = ~in[236]; 
    assign layer_0[1289] = ~(in[687] ^ in[795]); 
    assign layer_0[1290] = 1'b1; 
    assign layer_0[1291] = in[910] ^ in[70]; 
    assign layer_0[1292] = in[758] ^ in[570]; 
    assign layer_0[1293] = in[812] | in[696]; 
    assign layer_0[1294] = in[568] ^ in[94]; 
    assign layer_0[1295] = ~in[621] | (in[288] & in[621]); 
    assign layer_0[1296] = in[714] & ~in[478]; 
    assign layer_0[1297] = ~(in[934] ^ in[660]); 
    assign layer_0[1298] = ~(in[936] ^ in[583]); 
    assign layer_0[1299] = in[715] & in[583]; 
    assign layer_0[1300] = ~(in[276] & in[2]); 
    assign layer_0[1301] = in[5] ^ in[949]; 
    assign layer_0[1302] = in[1003] ^ in[381]; 
    assign layer_0[1303] = in[872]; 
    assign layer_0[1304] = ~in[25] | (in[939] & in[25]); 
    assign layer_0[1305] = in[587] & ~in[97]; 
    assign layer_0[1306] = in[535] ^ in[513]; 
    assign layer_0[1307] = ~in[904] | (in[904] & in[265]); 
    assign layer_0[1308] = ~in[89] | (in[387] & in[89]); 
    assign layer_0[1309] = ~(in[885] ^ in[612]); 
    assign layer_0[1310] = in[632]; 
    assign layer_0[1311] = in[966] | in[260]; 
    assign layer_0[1312] = ~(in[584] ^ in[793]); 
    assign layer_0[1313] = ~in[533]; 
    assign layer_0[1314] = ~(in[538] ^ in[477]); 
    assign layer_0[1315] = in[951] ^ in[332]; 
    assign layer_0[1316] = ~(in[506] | in[793]); 
    assign layer_0[1317] = in[505]; 
    assign layer_0[1318] = in[714]; 
    assign layer_0[1319] = in[903] ^ in[918]; 
    assign layer_0[1320] = in[612] ^ in[619]; 
    assign layer_0[1321] = in[380] & in[318]; 
    assign layer_0[1322] = ~in[371] | (in[817] & in[371]); 
    assign layer_0[1323] = in[145]; 
    assign layer_0[1324] = ~in[300]; 
    assign layer_0[1325] = in[31] ^ in[489]; 
    assign layer_0[1326] = in[246] ^ in[45]; 
    assign layer_0[1327] = ~in[265] | (in[265] & in[1013]); 
    assign layer_0[1328] = ~(in[551] ^ in[855]); 
    assign layer_0[1329] = in[345] & ~in[456]; 
    assign layer_0[1330] = in[534]; 
    assign layer_0[1331] = ~(in[600] ^ in[12]); 
    assign layer_0[1332] = ~in[577]; 
    assign layer_0[1333] = ~(in[600] ^ in[264]); 
    assign layer_0[1334] = in[634] ^ in[239]; 
    assign layer_0[1335] = in[689] ^ in[628]; 
    assign layer_0[1336] = in[479] | in[841]; 
    assign layer_0[1337] = in[776] | in[554]; 
    assign layer_0[1338] = ~in[986] | (in[382] & in[986]); 
    assign layer_0[1339] = in[1016] | in[491]; 
    assign layer_0[1340] = ~in[778]; 
    assign layer_0[1341] = ~in[632] | (in[493] & in[632]); 
    assign layer_0[1342] = ~(in[553] ^ in[46]); 
    assign layer_0[1343] = ~in[179] | (in[595] & in[179]); 
    assign layer_0[1344] = in[653] & ~in[901]; 
    assign layer_0[1345] = ~in[682]; 
    assign layer_0[1346] = in[809]; 
    assign layer_0[1347] = ~(in[478] | in[856]); 
    assign layer_0[1348] = ~in[340] | (in[87] & in[340]); 
    assign layer_0[1349] = ~in[611] | (in[989] & in[611]); 
    assign layer_0[1350] = in[541]; 
    assign layer_0[1351] = ~(in[619] ^ in[819]); 
    assign layer_0[1352] = in[647] & ~in[17]; 
    assign layer_0[1353] = ~in[9] | (in[954] & in[9]); 
    assign layer_0[1354] = in[675] & ~in[923]; 
    assign layer_0[1355] = in[103] & ~in[156]; 
    assign layer_0[1356] = in[743]; 
    assign layer_0[1357] = in[24] ^ in[1001]; 
    assign layer_0[1358] = in[165] ^ in[308]; 
    assign layer_0[1359] = in[730]; 
    assign layer_0[1360] = in[446] | in[1014]; 
    assign layer_0[1361] = in[573] ^ in[951]; 
    assign layer_0[1362] = ~(in[776] ^ in[1000]); 
    assign layer_0[1363] = in[951] ^ in[873]; 
    assign layer_0[1364] = in[764] & in[405]; 
    assign layer_0[1365] = in[407] & in[808]; 
    assign layer_0[1366] = in[537] ^ in[923]; 
    assign layer_0[1367] = in[666] ^ in[536]; 
    assign layer_0[1368] = in[564]; 
    assign layer_0[1369] = ~(in[330] ^ in[632]); 
    assign layer_0[1370] = ~in[321]; 
    assign layer_0[1371] = in[740]; 
    assign layer_0[1372] = in[389] & in[838]; 
    assign layer_0[1373] = ~(in[474] | in[988]); 
    assign layer_0[1374] = ~in[741]; 
    assign layer_0[1375] = in[405] & ~in[191]; 
    assign layer_0[1376] = ~(in[206] ^ in[700]); 
    assign layer_0[1377] = ~(in[687] & in[134]); 
    assign layer_0[1378] = ~in[792] | (in[699] & in[792]); 
    assign layer_0[1379] = in[558] | in[611]; 
    assign layer_0[1380] = in[729] & ~in[532]; 
    assign layer_0[1381] = in[393]; 
    assign layer_0[1382] = ~(in[47] & in[422]); 
    assign layer_0[1383] = in[402] | in[78]; 
    assign layer_0[1384] = in[414] ^ in[664]; 
    assign layer_0[1385] = in[830] & ~in[273]; 
    assign layer_0[1386] = in[677] ^ in[264]; 
    assign layer_0[1387] = in[824] ^ in[875]; 
    assign layer_0[1388] = in[991] & in[342]; 
    assign layer_0[1389] = ~(in[385] ^ in[805]); 
    assign layer_0[1390] = ~in[724] | (in[222] & in[724]); 
    assign layer_0[1391] = in[824] & in[264]; 
    assign layer_0[1392] = in[592]; 
    assign layer_0[1393] = in[205] ^ in[892]; 
    assign layer_0[1394] = ~(in[590] | in[99]); 
    assign layer_0[1395] = in[347]; 
    assign layer_0[1396] = in[299] ^ in[552]; 
    assign layer_0[1397] = ~(in[990] ^ in[933]); 
    assign layer_0[1398] = in[731] ^ in[980]; 
    assign layer_0[1399] = in[869] | in[49]; 
    assign layer_0[1400] = ~(in[1022] | in[251]); 
    assign layer_0[1401] = ~in[950]; 
    assign layer_0[1402] = ~(in[597] & in[730]); 
    assign layer_0[1403] = ~(in[472] ^ in[930]); 
    assign layer_0[1404] = in[178] ^ in[441]; 
    assign layer_0[1405] = in[745] ^ in[711]; 
    assign layer_0[1406] = ~(in[113] ^ in[519]); 
    assign layer_0[1407] = ~(in[751] | in[518]); 
    assign layer_0[1408] = in[588] ^ in[969]; 
    assign layer_0[1409] = ~in[792]; 
    assign layer_0[1410] = ~(in[877] & in[93]); 
    assign layer_0[1411] = ~in[640] | (in[640] & in[1007]); 
    assign layer_0[1412] = in[222] ^ in[697]; 
    assign layer_0[1413] = ~(in[225] ^ in[457]); 
    assign layer_0[1414] = ~(in[163] & in[234]); 
    assign layer_0[1415] = in[610] ^ in[331]; 
    assign layer_0[1416] = in[413] | in[980]; 
    assign layer_0[1417] = ~(in[666] ^ in[285]); 
    assign layer_0[1418] = in[875] | in[656]; 
    assign layer_0[1419] = in[709] ^ in[759]; 
    assign layer_0[1420] = ~(in[520] ^ in[291]); 
    assign layer_0[1421] = ~in[508] | (in[508] & in[505]); 
    assign layer_0[1422] = ~(in[488] & in[455]); 
    assign layer_0[1423] = in[132] ^ in[6]; 
    assign layer_0[1424] = in[309] | in[11]; 
    assign layer_0[1425] = ~in[62] | (in[62] & in[991]); 
    assign layer_0[1426] = in[558]; 
    assign layer_0[1427] = in[829]; 
    assign layer_0[1428] = ~(in[588] ^ in[925]); 
    assign layer_0[1429] = in[634] ^ in[493]; 
    assign layer_0[1430] = in[358] ^ in[354]; 
    assign layer_0[1431] = in[160] & ~in[611]; 
    assign layer_0[1432] = ~(in[598] ^ in[584]); 
    assign layer_0[1433] = in[263] & ~in[300]; 
    assign layer_0[1434] = ~(in[480] & in[304]); 
    assign layer_0[1435] = ~(in[708] ^ in[546]); 
    assign layer_0[1436] = in[586] & in[586]; 
    assign layer_0[1437] = 1'b0; 
    assign layer_0[1438] = in[333] & ~in[129]; 
    assign layer_0[1439] = in[774] | in[82]; 
    assign layer_0[1440] = in[965]; 
    assign layer_0[1441] = in[316] | in[658]; 
    assign layer_0[1442] = ~in[387]; 
    assign layer_0[1443] = ~(in[768] | in[691]); 
    assign layer_0[1444] = in[259] ^ in[618]; 
    assign layer_0[1445] = in[764] ^ in[208]; 
    assign layer_0[1446] = ~in[712] | (in[461] & in[712]); 
    assign layer_0[1447] = in[458]; 
    assign layer_0[1448] = in[853] & ~in[640]; 
    assign layer_0[1449] = in[295] & ~in[1016]; 
    assign layer_0[1450] = ~in[180] | (in[715] & in[180]); 
    assign layer_0[1451] = in[800] & in[396]; 
    assign layer_0[1452] = ~in[412] | (in[412] & in[1018]); 
    assign layer_0[1453] = ~in[810]; 
    assign layer_0[1454] = ~(in[161] ^ in[678]); 
    assign layer_0[1455] = ~in[674]; 
    assign layer_0[1456] = 1'b0; 
    assign layer_0[1457] = ~in[209]; 
    assign layer_0[1458] = ~(in[1017] ^ in[1001]); 
    assign layer_0[1459] = in[371] & ~in[660]; 
    assign layer_0[1460] = ~(in[777] ^ in[755]); 
    assign layer_0[1461] = ~(in[891] | in[886]); 
    assign layer_0[1462] = ~(in[588] | in[557]); 
    assign layer_0[1463] = in[286]; 
    assign layer_0[1464] = ~(in[819] ^ in[499]); 
    assign layer_0[1465] = in[663]; 
    assign layer_0[1466] = ~(in[885] ^ in[127]); 
    assign layer_0[1467] = in[246]; 
    assign layer_0[1468] = in[197] & in[860]; 
    assign layer_0[1469] = in[946] | in[365]; 
    assign layer_0[1470] = ~(in[999] ^ in[379]); 
    assign layer_0[1471] = ~in[397]; 
    assign layer_0[1472] = ~in[666] | (in[666] & in[596]); 
    assign layer_0[1473] = ~in[58] | (in[58] & in[84]); 
    assign layer_0[1474] = in[649] & in[282]; 
    assign layer_0[1475] = in[820] ^ in[804]; 
    assign layer_0[1476] = in[429] ^ in[772]; 
    assign layer_0[1477] = ~(in[350] | in[226]); 
    assign layer_0[1478] = in[296] & ~in[307]; 
    assign layer_0[1479] = ~in[517]; 
    assign layer_0[1480] = ~in[216] | (in[667] & in[216]); 
    assign layer_0[1481] = in[326] & ~in[769]; 
    assign layer_0[1482] = in[765]; 
    assign layer_0[1483] = in[926] & ~in[69]; 
    assign layer_0[1484] = ~(in[177] | in[1010]); 
    assign layer_0[1485] = ~in[692]; 
    assign layer_0[1486] = ~(in[348] & in[284]); 
    assign layer_0[1487] = ~in[763]; 
    assign layer_0[1488] = in[395] & ~in[803]; 
    assign layer_0[1489] = in[598] ^ in[455]; 
    assign layer_0[1490] = ~(in[108] ^ in[214]); 
    assign layer_0[1491] = ~(in[533] ^ in[792]); 
    assign layer_0[1492] = ~(in[916] ^ in[279]); 
    assign layer_0[1493] = ~(in[662] & in[19]); 
    assign layer_0[1494] = ~(in[296] & in[333]); 
    assign layer_0[1495] = 1'b1; 
    assign layer_0[1496] = ~(in[857] ^ in[1015]); 
    assign layer_0[1497] = ~(in[499] | in[508]); 
    assign layer_0[1498] = ~(in[922] | in[709]); 
    assign layer_0[1499] = in[834] ^ in[340]; 
    assign layer_0[1500] = in[949] ^ in[936]; 
    assign layer_0[1501] = ~(in[985] | in[130]); 
    assign layer_0[1502] = in[63] | in[384]; 
    assign layer_0[1503] = in[66] & in[613]; 
    assign layer_0[1504] = ~(in[587] ^ in[667]); 
    assign layer_0[1505] = in[606] ^ in[196]; 
    assign layer_0[1506] = in[205] & ~in[977]; 
    assign layer_0[1507] = ~in[710] | (in[710] & in[681]); 
    assign layer_0[1508] = ~in[986] | (in[691] & in[986]); 
    assign layer_0[1509] = in[232] & ~in[965]; 
    assign layer_0[1510] = in[46] & ~in[536]; 
    assign layer_0[1511] = ~(in[53] ^ in[428]); 
    assign layer_0[1512] = in[952] ^ in[521]; 
    assign layer_0[1513] = in[1005] | in[953]; 
    assign layer_0[1514] = ~in[778]; 
    assign layer_0[1515] = in[397] & in[82]; 
    assign layer_0[1516] = in[163] ^ in[34]; 
    assign layer_0[1517] = ~(in[1003] | in[65]); 
    assign layer_0[1518] = in[621] & in[439]; 
    assign layer_0[1519] = ~(in[930] ^ in[841]); 
    assign layer_0[1520] = ~(in[612] ^ in[180]); 
    assign layer_0[1521] = in[372] ^ in[965]; 
    assign layer_0[1522] = in[348]; 
    assign layer_0[1523] = ~in[325] | (in[325] & in[557]); 
    assign layer_0[1524] = ~(in[352] & in[916]); 
    assign layer_0[1525] = ~in[400]; 
    assign layer_0[1526] = ~(in[601] & in[600]); 
    assign layer_0[1527] = in[948] ^ in[434]; 
    assign layer_0[1528] = ~(in[669] ^ in[550]); 
    assign layer_0[1529] = in[209] & in[345]; 
    assign layer_0[1530] = in[94] & ~in[276]; 
    assign layer_0[1531] = in[519] ^ in[539]; 
    assign layer_0[1532] = ~in[679]; 
    assign layer_0[1533] = in[893] ^ in[291]; 
    assign layer_0[1534] = in[974] & in[228]; 
    assign layer_0[1535] = in[260] & in[326]; 
    assign layer_0[1536] = in[632] ^ in[633]; 
    assign layer_0[1537] = ~(in[853] ^ in[837]); 
    assign layer_0[1538] = ~in[570]; 
    assign layer_0[1539] = in[461]; 
    assign layer_0[1540] = ~(in[935] | in[977]); 
    assign layer_0[1541] = ~(in[882] ^ in[222]); 
    assign layer_0[1542] = in[806] & ~in[670]; 
    assign layer_0[1543] = in[653] & ~in[1011]; 
    assign layer_0[1544] = in[949] & in[399]; 
    assign layer_0[1545] = ~(in[907] ^ in[284]); 
    assign layer_0[1546] = ~(in[628] ^ in[530]); 
    assign layer_0[1547] = ~(in[537] ^ in[474]); 
    assign layer_0[1548] = ~in[386] | (in[386] & in[526]); 
    assign layer_0[1549] = in[7] ^ in[752]; 
    assign layer_0[1550] = ~in[886] | (in[1003] & in[886]); 
    assign layer_0[1551] = ~(in[1018] & in[265]); 
    assign layer_0[1552] = in[238] | in[876]; 
    assign layer_0[1553] = ~(in[907] ^ in[637]); 
    assign layer_0[1554] = ~(in[601] & in[937]); 
    assign layer_0[1555] = ~(in[793] | in[716]); 
    assign layer_0[1556] = in[292] & in[502]; 
    assign layer_0[1557] = ~in[699] | (in[324] & in[699]); 
    assign layer_0[1558] = ~in[595] | (in[910] & in[595]); 
    assign layer_0[1559] = ~(in[331] ^ in[840]); 
    assign layer_0[1560] = ~in[713] | (in[291] & in[713]); 
    assign layer_0[1561] = in[521] & ~in[776]; 
    assign layer_0[1562] = in[492] ^ in[747]; 
    assign layer_0[1563] = ~in[228] | (in[228] & in[18]); 
    assign layer_0[1564] = ~(in[983] ^ in[984]); 
    assign layer_0[1565] = ~(in[432] & in[772]); 
    assign layer_0[1566] = in[710] ^ in[490]; 
    assign layer_0[1567] = ~in[746] | (in[264] & in[746]); 
    assign layer_0[1568] = ~(in[862] ^ in[584]); 
    assign layer_0[1569] = ~in[540] | (in[703] & in[540]); 
    assign layer_0[1570] = ~in[44] | (in[801] & in[44]); 
    assign layer_0[1571] = in[851] & in[588]; 
    assign layer_0[1572] = in[516] & ~in[754]; 
    assign layer_0[1573] = ~in[823]; 
    assign layer_0[1574] = ~(in[252] & in[508]); 
    assign layer_0[1575] = in[1016]; 
    assign layer_0[1576] = in[445] ^ in[677]; 
    assign layer_0[1577] = in[413] & in[602]; 
    assign layer_0[1578] = ~in[125]; 
    assign layer_0[1579] = ~(in[134] ^ in[710]); 
    assign layer_0[1580] = ~in[673] | (in[673] & in[292]); 
    assign layer_0[1581] = ~in[859]; 
    assign layer_0[1582] = ~(in[617] ^ in[919]); 
    assign layer_0[1583] = ~(in[173] ^ in[459]); 
    assign layer_0[1584] = ~in[300] | (in[300] & in[841]); 
    assign layer_0[1585] = in[921] | in[776]; 
    assign layer_0[1586] = in[470] & ~in[492]; 
    assign layer_0[1587] = ~in[809] | (in[809] & in[707]); 
    assign layer_0[1588] = in[213] ^ in[573]; 
    assign layer_0[1589] = ~(in[654] ^ in[887]); 
    assign layer_0[1590] = in[151] & ~in[279]; 
    assign layer_0[1591] = ~in[748]; 
    assign layer_0[1592] = ~(in[872] | in[837]); 
    assign layer_0[1593] = in[743] & in[82]; 
    assign layer_0[1594] = ~(in[624] | in[728]); 
    assign layer_0[1595] = in[205] ^ in[689]; 
    assign layer_0[1596] = ~in[19]; 
    assign layer_0[1597] = in[999]; 
    assign layer_0[1598] = in[789] & in[693]; 
    assign layer_0[1599] = in[920] & ~in[789]; 
    assign layer_0[1600] = in[864] & ~in[554]; 
    assign layer_0[1601] = ~(in[329] | in[563]); 
    assign layer_0[1602] = in[330] ^ in[876]; 
    assign layer_0[1603] = in[761] & in[835]; 
    assign layer_0[1604] = in[503] | in[840]; 
    assign layer_0[1605] = ~(in[452] ^ in[756]); 
    assign layer_0[1606] = ~(in[909] | in[240]); 
    assign layer_0[1607] = ~in[19] | (in[529] & in[19]); 
    assign layer_0[1608] = ~in[827] | (in[403] & in[827]); 
    assign layer_0[1609] = in[161] & in[487]; 
    assign layer_0[1610] = in[893] & ~in[948]; 
    assign layer_0[1611] = ~(in[933] ^ in[580]); 
    assign layer_0[1612] = in[540] ^ in[873]; 
    assign layer_0[1613] = in[588] ^ in[700]; 
    assign layer_0[1614] = in[855] & ~in[256]; 
    assign layer_0[1615] = ~(in[374] & in[376]); 
    assign layer_0[1616] = ~(in[880] & in[933]); 
    assign layer_0[1617] = in[515] & ~in[1013]; 
    assign layer_0[1618] = in[283] & in[149]; 
    assign layer_0[1619] = in[909]; 
    assign layer_0[1620] = ~(in[94] ^ in[395]); 
    assign layer_0[1621] = ~in[932] | (in[268] & in[932]); 
    assign layer_0[1622] = ~(in[208] ^ in[316]); 
    assign layer_0[1623] = ~(in[905] | in[508]); 
    assign layer_0[1624] = in[737] & in[430]; 
    assign layer_0[1625] = in[886] ^ in[250]; 
    assign layer_0[1626] = ~in[50] | (in[317] & in[50]); 
    assign layer_0[1627] = in[839] & ~in[826]; 
    assign layer_0[1628] = in[733] & in[17]; 
    assign layer_0[1629] = in[725] ^ in[316]; 
    assign layer_0[1630] = ~in[635] | (in[253] & in[635]); 
    assign layer_0[1631] = ~in[438] | (in[28] & in[438]); 
    assign layer_0[1632] = ~(in[237] & in[412]); 
    assign layer_0[1633] = in[808] ^ in[806]; 
    assign layer_0[1634] = in[663] & ~in[480]; 
    assign layer_0[1635] = ~(in[204] | in[248]); 
    assign layer_0[1636] = ~(in[701] | in[322]); 
    assign layer_0[1637] = ~(in[0] | in[525]); 
    assign layer_0[1638] = ~(in[872] & in[839]); 
    assign layer_0[1639] = ~(in[650] ^ in[757]); 
    assign layer_0[1640] = ~(in[746] ^ in[34]); 
    assign layer_0[1641] = in[331] ^ in[209]; 
    assign layer_0[1642] = 1'b1; 
    assign layer_0[1643] = ~in[491] | (in[491] & in[973]); 
    assign layer_0[1644] = ~(in[948] ^ in[101]); 
    assign layer_0[1645] = in[195] ^ in[583]; 
    assign layer_0[1646] = ~(in[821] ^ in[474]); 
    assign layer_0[1647] = ~(in[941] ^ in[462]); 
    assign layer_0[1648] = ~in[707] | (in[98] & in[707]); 
    assign layer_0[1649] = in[685]; 
    assign layer_0[1650] = ~(in[690] | in[938]); 
    assign layer_0[1651] = in[290] ^ in[803]; 
    assign layer_0[1652] = ~(in[244] & in[130]); 
    assign layer_0[1653] = in[739] | in[980]; 
    assign layer_0[1654] = ~(in[527] ^ in[780]); 
    assign layer_0[1655] = 1'b0; 
    assign layer_0[1656] = ~(in[391] ^ in[301]); 
    assign layer_0[1657] = ~(in[229] | in[899]); 
    assign layer_0[1658] = ~in[740] | (in[513] & in[740]); 
    assign layer_0[1659] = ~in[382]; 
    assign layer_0[1660] = ~(in[776] | in[578]); 
    assign layer_0[1661] = in[973] | in[731]; 
    assign layer_0[1662] = in[97]; 
    assign layer_0[1663] = ~(in[798] ^ in[297]); 
    assign layer_0[1664] = in[917] & ~in[868]; 
    assign layer_0[1665] = in[56] ^ in[242]; 
    assign layer_0[1666] = ~(in[755] ^ in[899]); 
    assign layer_0[1667] = in[371] ^ in[598]; 
    assign layer_0[1668] = in[40] & ~in[861]; 
    assign layer_0[1669] = in[397] ^ in[699]; 
    assign layer_0[1670] = ~(in[743] ^ in[573]); 
    assign layer_0[1671] = in[404] | in[526]; 
    assign layer_0[1672] = ~in[485]; 
    assign layer_0[1673] = in[630] ^ in[365]; 
    assign layer_0[1674] = ~in[871]; 
    assign layer_0[1675] = in[1]; 
    assign layer_0[1676] = in[795] & ~in[771]; 
    assign layer_0[1677] = ~(in[124] ^ in[223]); 
    assign layer_0[1678] = in[300] ^ in[887]; 
    assign layer_0[1679] = in[261] ^ in[18]; 
    assign layer_0[1680] = in[312] | in[824]; 
    assign layer_0[1681] = ~(in[600] ^ in[873]); 
    assign layer_0[1682] = ~(in[485] & in[227]); 
    assign layer_0[1683] = ~(in[504] | in[858]); 
    assign layer_0[1684] = in[713] ^ in[366]; 
    assign layer_0[1685] = ~(in[594] | in[910]); 
    assign layer_0[1686] = in[42] & in[580]; 
    assign layer_0[1687] = ~(in[614] ^ in[448]); 
    assign layer_0[1688] = ~in[324]; 
    assign layer_0[1689] = ~(in[556] & in[487]); 
    assign layer_0[1690] = in[730] & in[733]; 
    assign layer_0[1691] = in[662] ^ in[892]; 
    assign layer_0[1692] = in[208]; 
    assign layer_0[1693] = in[682] & ~in[94]; 
    assign layer_0[1694] = in[589] | in[277]; 
    assign layer_0[1695] = ~(in[603] & in[582]); 
    assign layer_0[1696] = ~(in[600] ^ in[648]); 
    assign layer_0[1697] = ~(in[871] ^ in[538]); 
    assign layer_0[1698] = ~in[53] | (in[30] & in[53]); 
    assign layer_0[1699] = in[82] & ~in[525]; 
    assign layer_0[1700] = ~(in[988] ^ in[194]); 
    assign layer_0[1701] = ~(in[632] | in[922]); 
    assign layer_0[1702] = in[360] & ~in[1]; 
    assign layer_0[1703] = ~(in[684] ^ in[645]); 
    assign layer_0[1704] = in[726]; 
    assign layer_0[1705] = in[35] & in[867]; 
    assign layer_0[1706] = ~in[673]; 
    assign layer_0[1707] = ~in[857]; 
    assign layer_0[1708] = in[636] ^ in[346]; 
    assign layer_0[1709] = in[694] & in[875]; 
    assign layer_0[1710] = in[789] ^ in[634]; 
    assign layer_0[1711] = ~in[976] | (in[907] & in[976]); 
    assign layer_0[1712] = ~in[870] | (in[870] & in[903]); 
    assign layer_0[1713] = in[613]; 
    assign layer_0[1714] = in[572] & ~in[481]; 
    assign layer_0[1715] = ~(in[805] ^ in[859]); 
    assign layer_0[1716] = in[1015] ^ in[563]; 
    assign layer_0[1717] = ~(in[351] ^ in[254]); 
    assign layer_0[1718] = ~in[327]; 
    assign layer_0[1719] = ~(in[878] ^ in[929]); 
    assign layer_0[1720] = in[127] ^ in[636]; 
    assign layer_0[1721] = in[55] ^ in[221]; 
    assign layer_0[1722] = in[535] & in[5]; 
    assign layer_0[1723] = in[730] & ~in[566]; 
    assign layer_0[1724] = in[641]; 
    assign layer_0[1725] = in[999] ^ in[718]; 
    assign layer_0[1726] = ~(in[795] ^ in[517]); 
    assign layer_0[1727] = in[713] ^ in[859]; 
    assign layer_0[1728] = ~(in[953] & in[121]); 
    assign layer_0[1729] = in[736] ^ in[255]; 
    assign layer_0[1730] = ~in[99] | (in[99] & in[432]); 
    assign layer_0[1731] = ~(in[741] ^ in[169]); 
    assign layer_0[1732] = in[328]; 
    assign layer_0[1733] = in[816] | in[397]; 
    assign layer_0[1734] = in[253] & ~in[589]; 
    assign layer_0[1735] = in[455] & ~in[56]; 
    assign layer_0[1736] = ~(in[35] | in[490]); 
    assign layer_0[1737] = ~in[888]; 
    assign layer_0[1738] = in[741] | in[256]; 
    assign layer_0[1739] = ~(in[947] ^ in[807]); 
    assign layer_0[1740] = in[723] ^ in[930]; 
    assign layer_0[1741] = ~in[315] | (in[315] & in[732]); 
    assign layer_0[1742] = in[822] ^ in[804]; 
    assign layer_0[1743] = ~(in[896] ^ in[931]); 
    assign layer_0[1744] = in[865] ^ in[582]; 
    assign layer_0[1745] = in[300] | in[27]; 
    assign layer_0[1746] = ~(in[643] ^ in[283]); 
    assign layer_0[1747] = in[443]; 
    assign layer_0[1748] = ~in[888] | (in[640] & in[888]); 
    assign layer_0[1749] = in[577]; 
    assign layer_0[1750] = in[933] & ~in[763]; 
    assign layer_0[1751] = ~(in[318] & in[280]); 
    assign layer_0[1752] = in[567] ^ in[892]; 
    assign layer_0[1753] = in[806]; 
    assign layer_0[1754] = in[345] & ~in[552]; 
    assign layer_0[1755] = in[372] ^ in[612]; 
    assign layer_0[1756] = in[849] | in[322]; 
    assign layer_0[1757] = in[20] & ~in[652]; 
    assign layer_0[1758] = ~(in[654] | in[986]); 
    assign layer_0[1759] = ~(in[498] ^ in[516]); 
    assign layer_0[1760] = ~in[824]; 
    assign layer_0[1761] = ~(in[224] & in[292]); 
    assign layer_0[1762] = ~(in[29] | in[319]); 
    assign layer_0[1763] = in[920] ^ in[918]; 
    assign layer_0[1764] = in[653]; 
    assign layer_0[1765] = ~(in[1014] ^ in[923]); 
    assign layer_0[1766] = ~(in[688] ^ in[718]); 
    assign layer_0[1767] = in[919] ^ in[871]; 
    assign layer_0[1768] = ~(in[519] ^ in[97]); 
    assign layer_0[1769] = ~(in[809] ^ in[517]); 
    assign layer_0[1770] = in[860] | in[843]; 
    assign layer_0[1771] = in[499] | in[965]; 
    assign layer_0[1772] = in[298] & ~in[734]; 
    assign layer_0[1773] = ~(in[324] ^ in[897]); 
    assign layer_0[1774] = in[445] ^ in[846]; 
    assign layer_0[1775] = ~(in[822] ^ in[999]); 
    assign layer_0[1776] = ~in[127] | (in[1008] & in[127]); 
    assign layer_0[1777] = ~in[27]; 
    assign layer_0[1778] = ~in[285]; 
    assign layer_0[1779] = in[287] & ~in[606]; 
    assign layer_0[1780] = in[84] | in[222]; 
    assign layer_0[1781] = ~(in[98] ^ in[929]); 
    assign layer_0[1782] = in[841] ^ in[886]; 
    assign layer_0[1783] = in[776]; 
    assign layer_0[1784] = in[150] & in[903]; 
    assign layer_0[1785] = in[473] ^ in[438]; 
    assign layer_0[1786] = ~in[415] | (in[63] & in[415]); 
    assign layer_0[1787] = in[39]; 
    assign layer_0[1788] = in[824]; 
    assign layer_0[1789] = in[77] ^ in[647]; 
    assign layer_0[1790] = ~in[902] | (in[938] & in[902]); 
    assign layer_0[1791] = in[878] | in[531]; 
    assign layer_0[1792] = in[654]; 
    assign layer_0[1793] = in[698] ^ in[459]; 
    assign layer_0[1794] = ~(in[568] ^ in[600]); 
    assign layer_0[1795] = in[743] & ~in[268]; 
    assign layer_0[1796] = ~(in[729] ^ in[582]); 
    assign layer_0[1797] = in[332]; 
    assign layer_0[1798] = ~(in[720] & in[941]); 
    assign layer_0[1799] = ~(in[835] ^ in[416]); 
    assign layer_0[1800] = in[949] & in[698]; 
    assign layer_0[1801] = in[123] ^ in[738]; 
    assign layer_0[1802] = ~in[499] | (in[499] & in[886]); 
    assign layer_0[1803] = ~in[6]; 
    assign layer_0[1804] = in[263] ^ in[762]; 
    assign layer_0[1805] = in[454] & ~in[51]; 
    assign layer_0[1806] = in[221] ^ in[127]; 
    assign layer_0[1807] = in[89]; 
    assign layer_0[1808] = ~(in[22] ^ in[691]); 
    assign layer_0[1809] = in[109]; 
    assign layer_0[1810] = ~(in[455] & in[297]); 
    assign layer_0[1811] = ~in[458] | (in[907] & in[458]); 
    assign layer_0[1812] = ~in[871]; 
    assign layer_0[1813] = ~in[836]; 
    assign layer_0[1814] = in[448] ^ in[733]; 
    assign layer_0[1815] = in[31] ^ in[667]; 
    assign layer_0[1816] = ~in[265]; 
    assign layer_0[1817] = ~in[647]; 
    assign layer_0[1818] = ~(in[899] & in[828]); 
    assign layer_0[1819] = in[36] ^ in[791]; 
    assign layer_0[1820] = in[688] & ~in[998]; 
    assign layer_0[1821] = in[713] | in[995]; 
    assign layer_0[1822] = in[1009] & in[894]; 
    assign layer_0[1823] = ~(in[336] | in[228]); 
    assign layer_0[1824] = in[952] & in[781]; 
    assign layer_0[1825] = ~(in[114] & in[403]); 
    assign layer_0[1826] = in[381]; 
    assign layer_0[1827] = ~(in[873] ^ in[730]); 
    assign layer_0[1828] = ~(in[797] | in[614]); 
    assign layer_0[1829] = in[46] | in[612]; 
    assign layer_0[1830] = in[146] & ~in[956]; 
    assign layer_0[1831] = ~(in[381] ^ in[939]); 
    assign layer_0[1832] = ~(in[673] & in[119]); 
    assign layer_0[1833] = in[839] & ~in[439]; 
    assign layer_0[1834] = ~in[867]; 
    assign layer_0[1835] = in[641]; 
    assign layer_0[1836] = in[493] ^ in[980]; 
    assign layer_0[1837] = ~(in[913] ^ in[931]); 
    assign layer_0[1838] = ~(in[844] ^ in[253]); 
    assign layer_0[1839] = in[338]; 
    assign layer_0[1840] = in[85]; 
    assign layer_0[1841] = in[501] ^ in[850]; 
    assign layer_0[1842] = in[30] & ~in[401]; 
    assign layer_0[1843] = in[924] ^ in[872]; 
    assign layer_0[1844] = ~in[634]; 
    assign layer_0[1845] = in[797]; 
    assign layer_0[1846] = ~in[915]; 
    assign layer_0[1847] = ~in[175]; 
    assign layer_0[1848] = ~in[877]; 
    assign layer_0[1849] = ~(in[411] & in[1022]); 
    assign layer_0[1850] = in[216] ^ in[826]; 
    assign layer_0[1851] = in[574] ^ in[964]; 
    assign layer_0[1852] = in[875] & ~in[500]; 
    assign layer_0[1853] = ~(in[705] | in[342]); 
    assign layer_0[1854] = in[608] ^ in[505]; 
    assign layer_0[1855] = in[979] ^ in[764]; 
    assign layer_0[1856] = ~(in[684] ^ in[161]); 
    assign layer_0[1857] = in[643] & ~in[266]; 
    assign layer_0[1858] = ~in[603]; 
    assign layer_0[1859] = in[218] & in[208]; 
    assign layer_0[1860] = in[442] & ~in[699]; 
    assign layer_0[1861] = in[203] & in[692]; 
    assign layer_0[1862] = in[241] ^ in[747]; 
    assign layer_0[1863] = ~(in[82] & in[107]); 
    assign layer_0[1864] = in[133] & ~in[937]; 
    assign layer_0[1865] = ~(in[535] ^ in[189]); 
    assign layer_0[1866] = in[763]; 
    assign layer_0[1867] = in[445]; 
    assign layer_0[1868] = ~in[11]; 
    assign layer_0[1869] = ~in[137] | (in[137] & in[967]); 
    assign layer_0[1870] = in[58] & ~in[805]; 
    assign layer_0[1871] = ~(in[767] & in[298]); 
    assign layer_0[1872] = ~(in[887] ^ in[873]); 
    assign layer_0[1873] = ~in[455] | (in[455] & in[363]); 
    assign layer_0[1874] = ~(in[802] ^ in[933]); 
    assign layer_0[1875] = ~in[153] | (in[153] & in[980]); 
    assign layer_0[1876] = ~in[856]; 
    assign layer_0[1877] = in[891] ^ in[260]; 
    assign layer_0[1878] = 1'b1; 
    assign layer_0[1879] = in[62] & ~in[720]; 
    assign layer_0[1880] = ~in[664]; 
    assign layer_0[1881] = ~(in[754] ^ in[381]); 
    assign layer_0[1882] = ~(in[897] | in[979]); 
    assign layer_0[1883] = ~in[284] | (in[284] & in[775]); 
    assign layer_0[1884] = ~in[166] | (in[929] & in[166]); 
    assign layer_0[1885] = in[757] ^ in[116]; 
    assign layer_0[1886] = ~(in[770] | in[473]); 
    assign layer_0[1887] = in[39] & ~in[548]; 
    assign layer_0[1888] = in[811] & ~in[875]; 
    assign layer_0[1889] = ~(in[683] ^ in[397]); 
    assign layer_0[1890] = ~in[443] | (in[443] & in[348]); 
    assign layer_0[1891] = in[442] & in[961]; 
    assign layer_0[1892] = ~(in[488] ^ in[310]); 
    assign layer_0[1893] = in[731] & in[413]; 
    assign layer_0[1894] = ~in[428] | (in[428] & in[827]); 
    assign layer_0[1895] = in[10] | in[676]; 
    assign layer_0[1896] = ~(in[103] & in[968]); 
    assign layer_0[1897] = ~(in[535] ^ in[228]); 
    assign layer_0[1898] = ~in[684]; 
    assign layer_0[1899] = ~(in[868] | in[295]); 
    assign layer_0[1900] = ~(in[337] ^ in[434]); 
    assign layer_0[1901] = in[629] | in[805]; 
    assign layer_0[1902] = ~in[613]; 
    assign layer_0[1903] = in[803] ^ in[627]; 
    assign layer_0[1904] = in[951] | in[793]; 
    assign layer_0[1905] = ~(in[68] ^ in[551]); 
    assign layer_0[1906] = in[549] ^ in[970]; 
    assign layer_0[1907] = ~in[997] | (in[49] & in[997]); 
    assign layer_0[1908] = ~in[861]; 
    assign layer_0[1909] = ~in[916]; 
    assign layer_0[1910] = ~in[644] | (in[852] & in[644]); 
    assign layer_0[1911] = ~(in[874] ^ in[584]); 
    assign layer_0[1912] = ~in[748] | (in[543] & in[748]); 
    assign layer_0[1913] = in[442] ^ in[649]; 
    assign layer_0[1914] = ~in[20]; 
    assign layer_0[1915] = in[548] ^ in[866]; 
    assign layer_0[1916] = ~(in[324] ^ in[915]); 
    assign layer_0[1917] = ~in[944] | (in[288] & in[944]); 
    assign layer_0[1918] = in[930] | in[762]; 
    assign layer_0[1919] = ~in[819] | (in[819] & in[804]); 
    assign layer_0[1920] = in[238]; 
    assign layer_0[1921] = in[388] | in[562]; 
    assign layer_0[1922] = ~(in[190] ^ in[264]); 
    assign layer_0[1923] = ~in[604]; 
    assign layer_0[1924] = in[173] & ~in[23]; 
    assign layer_0[1925] = ~(in[325] & in[445]); 
    assign layer_0[1926] = in[943] | in[912]; 
    assign layer_0[1927] = in[468] ^ in[774]; 
    assign layer_0[1928] = ~in[902] | (in[902] & in[878]); 
    assign layer_0[1929] = in[724] ^ in[79]; 
    assign layer_0[1930] = ~(in[888] ^ in[699]); 
    assign layer_0[1931] = in[953] & ~in[370]; 
    assign layer_0[1932] = ~in[1016] | (in[1016] & in[877]); 
    assign layer_0[1933] = in[844] & ~in[253]; 
    assign layer_0[1934] = ~(in[485] ^ in[504]); 
    assign layer_0[1935] = in[553]; 
    assign layer_0[1936] = ~in[470]; 
    assign layer_0[1937] = ~(in[129] ^ in[667]); 
    assign layer_0[1938] = in[958] ^ in[469]; 
    assign layer_0[1939] = ~(in[885] ^ in[872]); 
    assign layer_0[1940] = ~(in[552] ^ in[584]); 
    assign layer_0[1941] = ~(in[767] & in[151]); 
    assign layer_0[1942] = ~in[120]; 
    assign layer_0[1943] = in[362] ^ in[416]; 
    assign layer_0[1944] = in[13] ^ in[789]; 
    assign layer_0[1945] = in[1003] ^ in[81]; 
    assign layer_0[1946] = ~(in[804] | in[981]); 
    assign layer_0[1947] = in[598] & in[629]; 
    assign layer_0[1948] = in[659]; 
    assign layer_0[1949] = in[923] & ~in[988]; 
    assign layer_0[1950] = ~(in[550] | in[951]); 
    assign layer_0[1951] = in[916] ^ in[161]; 
    assign layer_0[1952] = ~(in[10] & in[629]); 
    assign layer_0[1953] = in[29] | in[321]; 
    assign layer_0[1954] = ~(in[78] ^ in[65]); 
    assign layer_0[1955] = ~in[826] | (in[826] & in[689]); 
    assign layer_0[1956] = ~(in[989] | in[679]); 
    assign layer_0[1957] = ~(in[30] ^ in[56]); 
    assign layer_0[1958] = in[344] & in[8]; 
    assign layer_0[1959] = ~in[317] | (in[473] & in[317]); 
    assign layer_0[1960] = in[714] & ~in[947]; 
    assign layer_0[1961] = in[415] ^ in[205]; 
    assign layer_0[1962] = ~(in[470] ^ in[599]); 
    assign layer_0[1963] = in[939] ^ in[626]; 
    assign layer_0[1964] = ~in[264]; 
    assign layer_0[1965] = ~(in[112] | in[1003]); 
    assign layer_0[1966] = ~in[901]; 
    assign layer_0[1967] = ~in[198]; 
    assign layer_0[1968] = ~(in[845] ^ in[282]); 
    assign layer_0[1969] = ~in[672] | (in[1] & in[672]); 
    assign layer_0[1970] = in[633]; 
    assign layer_0[1971] = in[341]; 
    assign layer_0[1972] = ~(in[284] ^ in[276]); 
    assign layer_0[1973] = ~(in[791] ^ in[517]); 
    assign layer_0[1974] = ~(in[722] ^ in[338]); 
    assign layer_0[1975] = ~(in[95] ^ in[159]); 
    assign layer_0[1976] = 1'b1; 
    assign layer_0[1977] = ~(in[952] | in[765]); 
    assign layer_0[1978] = ~in[356]; 
    assign layer_0[1979] = ~(in[684] ^ in[485]); 
    assign layer_0[1980] = ~(in[179] ^ in[659]); 
    assign layer_0[1981] = ~in[660] | (in[575] & in[660]); 
    assign layer_0[1982] = in[967] ^ in[469]; 
    assign layer_0[1983] = ~(in[935] | in[443]); 
    assign layer_0[1984] = ~(in[585] & in[664]); 
    assign layer_0[1985] = ~(in[615] ^ in[810]); 
    assign layer_0[1986] = in[915] & ~in[314]; 
    assign layer_0[1987] = in[41] & in[855]; 
    assign layer_0[1988] = ~in[970]; 
    assign layer_0[1989] = 1'b0; 
    assign layer_0[1990] = in[781] | in[681]; 
    assign layer_0[1991] = ~in[714]; 
    assign layer_0[1992] = in[963] & ~in[273]; 
    assign layer_0[1993] = ~in[3] | (in[78] & in[3]); 
    assign layer_0[1994] = in[311] & in[33]; 
    assign layer_0[1995] = in[10] ^ in[640]; 
    assign layer_0[1996] = in[937] & ~in[619]; 
    assign layer_0[1997] = in[314] ^ in[435]; 
    assign layer_0[1998] = ~(in[515] ^ in[446]); 
    assign layer_0[1999] = in[713] ^ in[883]; 
    assign layer_0[2000] = in[415] | in[533]; 
    assign layer_0[2001] = ~in[294] | (in[294] & in[366]); 
    assign layer_0[2002] = in[755] & ~in[920]; 
    assign layer_0[2003] = in[194] & ~in[260]; 
    assign layer_0[2004] = ~in[822]; 
    assign layer_0[2005] = ~in[455] | (in[455] & in[571]); 
    assign layer_0[2006] = in[1000] & ~in[593]; 
    assign layer_0[2007] = 1'b0; 
    assign layer_0[2008] = in[41] & in[422]; 
    assign layer_0[2009] = ~in[335] | (in[335] & in[798]); 
    assign layer_0[2010] = ~(in[250] ^ in[241]); 
    assign layer_0[2011] = in[184] ^ in[715]; 
    assign layer_0[2012] = ~in[962] | (in[765] & in[962]); 
    assign layer_0[2013] = in[804] & in[954]; 
    assign layer_0[2014] = ~(in[550] & in[981]); 
    assign layer_0[2015] = ~in[740]; 
    assign layer_0[2016] = in[217] & ~in[570]; 
    assign layer_0[2017] = ~(in[327] ^ in[506]); 
    assign layer_0[2018] = in[875] ^ in[730]; 
    assign layer_0[2019] = ~in[141] | (in[141] & in[916]); 
    assign layer_0[2020] = in[230] & ~in[327]; 
    assign layer_0[2021] = in[701]; 
    assign layer_0[2022] = in[642] & ~in[876]; 
    assign layer_0[2023] = in[324]; 
    assign layer_0[2024] = ~(in[629] ^ in[347]); 
    assign layer_0[2025] = ~in[177]; 
    assign layer_0[2026] = ~(in[951] ^ in[878]); 
    assign layer_0[2027] = ~in[1017] | (in[186] & in[1017]); 
    assign layer_0[2028] = ~(in[451] | in[668]); 
    assign layer_0[2029] = in[88] & in[184]; 
    assign layer_0[2030] = ~(in[709] ^ in[822]); 
    assign layer_0[2031] = in[996] | in[32]; 
    assign layer_0[2032] = in[940] ^ in[40]; 
    assign layer_0[2033] = in[821] | in[953]; 
    assign layer_0[2034] = ~(in[945] ^ in[652]); 
    assign layer_0[2035] = ~(in[939] ^ in[948]); 
    assign layer_0[2036] = in[762] ^ in[996]; 
    assign layer_0[2037] = in[236] ^ in[633]; 
    assign layer_0[2038] = ~(in[924] ^ in[13]); 
    assign layer_0[2039] = ~(in[920] ^ in[504]); 
    assign layer_0[2040] = in[146] & in[78]; 
    assign layer_0[2041] = in[232] & ~in[10]; 
    assign layer_0[2042] = ~in[38]; 
    assign layer_0[2043] = in[29]; 
    assign layer_0[2044] = ~(in[4] | in[504]); 
    assign layer_0[2045] = in[142] & in[661]; 
    assign layer_0[2046] = ~in[256]; 
    assign layer_0[2047] = ~(in[142] ^ in[759]); 
    assign layer_0[2048] = ~in[888]; 
    assign layer_0[2049] = ~(in[943] ^ in[717]); 
    assign layer_0[2050] = in[953] ^ in[98]; 
    assign layer_0[2051] = in[380] & ~in[159]; 
    assign layer_0[2052] = in[18] | in[825]; 
    assign layer_0[2053] = in[807]; 
    assign layer_0[2054] = in[970]; 
    assign layer_0[2055] = in[451] ^ in[322]; 
    assign layer_0[2056] = in[8] & in[427]; 
    assign layer_0[2057] = ~(in[905] ^ in[887]); 
    assign layer_0[2058] = in[1009] ^ in[97]; 
    assign layer_0[2059] = ~in[534]; 
    assign layer_0[2060] = ~(in[163] | in[419]); 
    assign layer_0[2061] = in[204]; 
    assign layer_0[2062] = in[364] & in[651]; 
    assign layer_0[2063] = ~in[664]; 
    assign layer_0[2064] = ~(in[8] ^ in[272]); 
    assign layer_0[2065] = in[355] ^ in[699]; 
    assign layer_0[2066] = in[398] & ~in[791]; 
    assign layer_0[2067] = in[668] | in[209]; 
    assign layer_0[2068] = in[449] ^ in[481]; 
    assign layer_0[2069] = in[896] | in[846]; 
    assign layer_0[2070] = ~(in[507] ^ in[429]); 
    assign layer_0[2071] = ~(in[905] ^ in[904]); 
    assign layer_0[2072] = in[900]; 
    assign layer_0[2073] = in[846]; 
    assign layer_0[2074] = ~(in[791] & in[1016]); 
    assign layer_0[2075] = in[560] & in[790]; 
    assign layer_0[2076] = 1'b0; 
    assign layer_0[2077] = in[979] | in[953]; 
    assign layer_0[2078] = in[913] | in[493]; 
    assign layer_0[2079] = ~in[478] | (in[46] & in[478]); 
    assign layer_0[2080] = in[547] & ~in[699]; 
    assign layer_0[2081] = in[996] & ~in[30]; 
    assign layer_0[2082] = in[597]; 
    assign layer_0[2083] = in[974] & in[913]; 
    assign layer_0[2084] = in[950] | in[1016]; 
    assign layer_0[2085] = in[728]; 
    assign layer_0[2086] = in[366] ^ in[266]; 
    assign layer_0[2087] = ~(in[953] ^ in[987]); 
    assign layer_0[2088] = in[445] ^ in[8]; 
    assign layer_0[2089] = ~in[376] | (in[795] & in[376]); 
    assign layer_0[2090] = ~(in[594] ^ in[888]); 
    assign layer_0[2091] = in[996] & in[236]; 
    assign layer_0[2092] = ~in[934] | (in[934] & in[62]); 
    assign layer_0[2093] = in[323] & ~in[29]; 
    assign layer_0[2094] = in[960] | in[38]; 
    assign layer_0[2095] = ~in[365] | (in[365] & in[837]); 
    assign layer_0[2096] = ~(in[612] | in[627]); 
    assign layer_0[2097] = ~(in[986] ^ in[985]); 
    assign layer_0[2098] = ~in[934] | (in[934] & in[935]); 
    assign layer_0[2099] = in[731]; 
    assign layer_0[2100] = in[825] ^ in[455]; 
    assign layer_0[2101] = ~in[840] | (in[184] & in[840]); 
    assign layer_0[2102] = in[623] & in[91]; 
    assign layer_0[2103] = ~(in[45] & in[338]); 
    assign layer_0[2104] = in[747] & in[381]; 
    assign layer_0[2105] = in[422] & ~in[1016]; 
    assign layer_0[2106] = in[648] ^ in[395]; 
    assign layer_0[2107] = in[856]; 
    assign layer_0[2108] = in[112]; 
    assign layer_0[2109] = ~(in[1017] ^ in[1016]); 
    assign layer_0[2110] = ~(in[970] ^ in[603]); 
    assign layer_0[2111] = in[217]; 
    assign layer_0[2112] = in[57] ^ in[957]; 
    assign layer_0[2113] = in[997] ^ in[18]; 
    assign layer_0[2114] = ~(in[279] ^ in[13]); 
    assign layer_0[2115] = ~in[889]; 
    assign layer_0[2116] = in[389] | in[618]; 
    assign layer_0[2117] = ~in[542] | (in[542] & in[625]); 
    assign layer_0[2118] = ~in[774]; 
    assign layer_0[2119] = in[519] & in[291]; 
    assign layer_0[2120] = ~(in[671] | in[840]); 
    assign layer_0[2121] = in[160] ^ in[263]; 
    assign layer_0[2122] = in[609] | in[693]; 
    assign layer_0[2123] = ~in[228] | (in[480] & in[228]); 
    assign layer_0[2124] = ~(in[926] ^ in[311]); 
    assign layer_0[2125] = 1'b0; 
    assign layer_0[2126] = ~(in[741] & in[791]); 
    assign layer_0[2127] = ~in[253] | (in[207] & in[253]); 
    assign layer_0[2128] = ~in[716] | (in[716] & in[322]); 
    assign layer_0[2129] = ~(in[49] ^ in[8]); 
    assign layer_0[2130] = ~(in[925] ^ in[590]); 
    assign layer_0[2131] = ~(in[253] | in[706]); 
    assign layer_0[2132] = in[825] ^ in[889]; 
    assign layer_0[2133] = ~(in[955] ^ in[692]); 
    assign layer_0[2134] = in[176] & in[339]; 
    assign layer_0[2135] = ~in[783] | (in[783] & in[274]); 
    assign layer_0[2136] = in[698] | in[6]; 
    assign layer_0[2137] = ~in[10] | (in[981] & in[10]); 
    assign layer_0[2138] = in[869] ^ in[254]; 
    assign layer_0[2139] = in[145] | in[577]; 
    assign layer_0[2140] = in[869] ^ in[67]; 
    assign layer_0[2141] = ~(in[609] ^ in[143]); 
    assign layer_0[2142] = ~(in[349] | in[332]); 
    assign layer_0[2143] = ~in[852]; 
    assign layer_0[2144] = in[1015]; 
    assign layer_0[2145] = in[662] & in[665]; 
    assign layer_0[2146] = ~(in[459] & in[359]); 
    assign layer_0[2147] = ~(in[582] ^ in[584]); 
    assign layer_0[2148] = in[52] ^ in[792]; 
    assign layer_0[2149] = in[822] | in[82]; 
    assign layer_0[2150] = ~(in[310] & in[653]); 
    assign layer_0[2151] = ~(in[266] & in[445]); 
    assign layer_0[2152] = in[984] & in[244]; 
    assign layer_0[2153] = ~(in[464] ^ in[460]); 
    assign layer_0[2154] = in[967]; 
    assign layer_0[2155] = in[969] ^ in[733]; 
    assign layer_0[2156] = in[492] & ~in[519]; 
    assign layer_0[2157] = ~in[387]; 
    assign layer_0[2158] = in[739] | in[315]; 
    assign layer_0[2159] = ~(in[932] | in[945]); 
    assign layer_0[2160] = ~(in[338] ^ in[959]); 
    assign layer_0[2161] = in[897]; 
    assign layer_0[2162] = in[299] & ~in[500]; 
    assign layer_0[2163] = in[768] | in[595]; 
    assign layer_0[2164] = ~(in[619] ^ in[708]); 
    assign layer_0[2165] = in[764] & in[666]; 
    assign layer_0[2166] = in[873] & ~in[954]; 
    assign layer_0[2167] = ~in[483] | (in[671] & in[483]); 
    assign layer_0[2168] = in[554] & ~in[364]; 
    assign layer_0[2169] = 1'b1; 
    assign layer_0[2170] = in[743] ^ in[261]; 
    assign layer_0[2171] = in[580] & ~in[762]; 
    assign layer_0[2172] = ~(in[334] & in[623]); 
    assign layer_0[2173] = 1'b0; 
    assign layer_0[2174] = ~(in[53] | in[232]); 
    assign layer_0[2175] = ~(in[931] ^ in[316]); 
    assign layer_0[2176] = in[349] ^ in[45]; 
    assign layer_0[2177] = in[931] | in[930]; 
    assign layer_0[2178] = in[68]; 
    assign layer_0[2179] = ~in[277] | (in[249] & in[277]); 
    assign layer_0[2180] = in[310] & in[850]; 
    assign layer_0[2181] = ~in[692]; 
    assign layer_0[2182] = ~(in[667] & in[402]); 
    assign layer_0[2183] = ~(in[626] ^ in[888]); 
    assign layer_0[2184] = in[96] | in[301]; 
    assign layer_0[2185] = ~in[954] | (in[692] & in[954]); 
    assign layer_0[2186] = ~in[505]; 
    assign layer_0[2187] = ~in[578]; 
    assign layer_0[2188] = in[266] | in[568]; 
    assign layer_0[2189] = ~(in[268] | in[966]); 
    assign layer_0[2190] = in[921]; 
    assign layer_0[2191] = ~(in[942] & in[643]); 
    assign layer_0[2192] = in[430]; 
    assign layer_0[2193] = ~(in[691] ^ in[749]); 
    assign layer_0[2194] = ~(in[574] | in[854]); 
    assign layer_0[2195] = in[268]; 
    assign layer_0[2196] = in[984] & ~in[833]; 
    assign layer_0[2197] = in[181] & in[509]; 
    assign layer_0[2198] = in[269] | in[144]; 
    assign layer_0[2199] = in[490] | in[882]; 
    assign layer_0[2200] = in[246] & ~in[792]; 
    assign layer_0[2201] = in[878] | in[20]; 
    assign layer_0[2202] = in[926] ^ in[590]; 
    assign layer_0[2203] = 1'b0; 
    assign layer_0[2204] = in[647] & ~in[624]; 
    assign layer_0[2205] = in[370] ^ in[569]; 
    assign layer_0[2206] = ~(in[682] ^ in[236]); 
    assign layer_0[2207] = in[780] ^ in[738]; 
    assign layer_0[2208] = in[508] ^ in[509]; 
    assign layer_0[2209] = 1'b1; 
    assign layer_0[2210] = in[448] & ~in[848]; 
    assign layer_0[2211] = in[23] ^ in[404]; 
    assign layer_0[2212] = ~(in[380] & in[972]); 
    assign layer_0[2213] = ~(in[870] ^ in[808]); 
    assign layer_0[2214] = in[1016] ^ in[921]; 
    assign layer_0[2215] = ~(in[824] ^ in[836]); 
    assign layer_0[2216] = ~in[197]; 
    assign layer_0[2217] = in[865] & ~in[653]; 
    assign layer_0[2218] = ~in[591] | (in[747] & in[591]); 
    assign layer_0[2219] = ~(in[984] ^ in[985]); 
    assign layer_0[2220] = ~in[969] | (in[287] & in[969]); 
    assign layer_0[2221] = ~(in[460] ^ in[712]); 
    assign layer_0[2222] = in[193]; 
    assign layer_0[2223] = ~(in[894] & in[958]); 
    assign layer_0[2224] = in[548] & ~in[948]; 
    assign layer_0[2225] = in[826] ^ in[985]; 
    assign layer_0[2226] = ~(in[265] ^ in[326]); 
    assign layer_0[2227] = ~in[25] | (in[771] & in[25]); 
    assign layer_0[2228] = ~in[324] | (in[882] & in[324]); 
    assign layer_0[2229] = ~(in[219] & in[476]); 
    assign layer_0[2230] = in[1001] ^ in[967]; 
    assign layer_0[2231] = in[514] | in[1012]; 
    assign layer_0[2232] = ~(in[765] ^ in[764]); 
    assign layer_0[2233] = in[27]; 
    assign layer_0[2234] = ~(in[625] ^ in[588]); 
    assign layer_0[2235] = in[110] & ~in[708]; 
    assign layer_0[2236] = in[661] & ~in[29]; 
    assign layer_0[2237] = in[346]; 
    assign layer_0[2238] = ~(in[359] & in[123]); 
    assign layer_0[2239] = in[181] & in[623]; 
    assign layer_0[2240] = in[587] & ~in[435]; 
    assign layer_0[2241] = ~(in[856] | in[856]); 
    assign layer_0[2242] = in[507] ^ in[148]; 
    assign layer_0[2243] = in[243] ^ in[848]; 
    assign layer_0[2244] = ~(in[208] ^ in[385]); 
    assign layer_0[2245] = ~in[263] | (in[3] & in[263]); 
    assign layer_0[2246] = in[345] & in[118]; 
    assign layer_0[2247] = ~(in[589] & in[323]); 
    assign layer_0[2248] = in[252]; 
    assign layer_0[2249] = in[507] | in[337]; 
    assign layer_0[2250] = ~(in[851] ^ in[195]); 
    assign layer_0[2251] = in[823] | in[402]; 
    assign layer_0[2252] = ~in[383] | (in[4] & in[383]); 
    assign layer_0[2253] = ~in[627]; 
    assign layer_0[2254] = in[360] ^ in[299]; 
    assign layer_0[2255] = in[696] ^ in[967]; 
    assign layer_0[2256] = ~(in[364] & in[260]); 
    assign layer_0[2257] = ~(in[246] ^ in[583]); 
    assign layer_0[2258] = ~in[166] | (in[166] & in[638]); 
    assign layer_0[2259] = in[977] | in[217]; 
    assign layer_0[2260] = in[4]; 
    assign layer_0[2261] = 1'b0; 
    assign layer_0[2262] = in[46] | in[337]; 
    assign layer_0[2263] = ~(in[953] ^ in[253]); 
    assign layer_0[2264] = ~(in[759] ^ in[603]); 
    assign layer_0[2265] = ~(in[265] & in[937]); 
    assign layer_0[2266] = in[115] ^ in[492]; 
    assign layer_0[2267] = ~in[327] | (in[327] & in[836]); 
    assign layer_0[2268] = in[827]; 
    assign layer_0[2269] = ~in[137] | (in[137] & in[716]); 
    assign layer_0[2270] = in[616] ^ in[637]; 
    assign layer_0[2271] = ~(in[234] ^ in[354]); 
    assign layer_0[2272] = ~(in[495] ^ in[39]); 
    assign layer_0[2273] = ~in[173]; 
    assign layer_0[2274] = in[907] ^ in[711]; 
    assign layer_0[2275] = ~(in[712] & in[157]); 
    assign layer_0[2276] = ~(in[1003] & in[519]); 
    assign layer_0[2277] = in[1008] & ~in[761]; 
    assign layer_0[2278] = ~(in[670] | in[872]); 
    assign layer_0[2279] = in[100] & ~in[33]; 
    assign layer_0[2280] = ~(in[997] ^ in[653]); 
    assign layer_0[2281] = ~in[347] | (in[347] & in[765]); 
    assign layer_0[2282] = in[627] ^ in[549]; 
    assign layer_0[2283] = ~in[437] | (in[211] & in[437]); 
    assign layer_0[2284] = in[355] & ~in[530]; 
    assign layer_0[2285] = in[340] & in[597]; 
    assign layer_0[2286] = in[242] ^ in[936]; 
    assign layer_0[2287] = in[969] & ~in[764]; 
    assign layer_0[2288] = in[467]; 
    assign layer_0[2289] = ~(in[911] ^ in[499]); 
    assign layer_0[2290] = ~(in[756] | in[125]); 
    assign layer_0[2291] = in[477] | in[825]; 
    assign layer_0[2292] = ~in[924]; 
    assign layer_0[2293] = in[522] | in[480]; 
    assign layer_0[2294] = in[266] & ~in[311]; 
    assign layer_0[2295] = in[798] ^ in[939]; 
    assign layer_0[2296] = in[35] & in[451]; 
    assign layer_0[2297] = in[808] ^ in[789]; 
    assign layer_0[2298] = in[90] ^ in[5]; 
    assign layer_0[2299] = in[393] & ~in[724]; 
    assign layer_0[2300] = in[480] & ~in[603]; 
    assign layer_0[2301] = ~(in[953] ^ in[555]); 
    assign layer_0[2302] = ~in[904]; 
    assign layer_0[2303] = ~(in[889] ^ in[715]); 
    assign layer_0[2304] = ~(in[162] ^ in[874]); 
    assign layer_0[2305] = ~in[977] | (in[461] & in[977]); 
    assign layer_0[2306] = in[765] ^ in[741]; 
    assign layer_0[2307] = ~in[950]; 
    assign layer_0[2308] = ~(in[864] ^ in[104]); 
    assign layer_0[2309] = in[343] & ~in[837]; 
    assign layer_0[2310] = in[69] ^ in[234]; 
    assign layer_0[2311] = in[986] ^ in[728]; 
    assign layer_0[2312] = ~(in[109] ^ in[1015]); 
    assign layer_0[2313] = in[1014] ^ in[397]; 
    assign layer_0[2314] = in[857] | in[985]; 
    assign layer_0[2315] = ~(in[309] | in[730]); 
    assign layer_0[2316] = ~in[557] | (in[557] & in[285]); 
    assign layer_0[2317] = ~in[401] | (in[401] & in[614]); 
    assign layer_0[2318] = ~in[484] | (in[765] & in[484]); 
    assign layer_0[2319] = in[60] ^ in[870]; 
    assign layer_0[2320] = ~in[536] | (in[536] & in[588]); 
    assign layer_0[2321] = ~in[535] | (in[535] & in[752]); 
    assign layer_0[2322] = ~(in[917] | in[777]); 
    assign layer_0[2323] = in[639] | in[484]; 
    assign layer_0[2324] = ~in[30]; 
    assign layer_0[2325] = in[264] & in[268]; 
    assign layer_0[2326] = ~in[962] | (in[962] & in[235]); 
    assign layer_0[2327] = ~(in[20] | in[533]); 
    assign layer_0[2328] = ~(in[600] & in[669]); 
    assign layer_0[2329] = in[385]; 
    assign layer_0[2330] = ~(in[40] | in[251]); 
    assign layer_0[2331] = in[457] & in[367]; 
    assign layer_0[2332] = ~in[605]; 
    assign layer_0[2333] = in[473] & ~in[100]; 
    assign layer_0[2334] = in[311] ^ in[478]; 
    assign layer_0[2335] = in[555] ^ in[520]; 
    assign layer_0[2336] = in[385] ^ in[175]; 
    assign layer_0[2337] = ~(in[971] ^ in[623]); 
    assign layer_0[2338] = in[259] ^ in[207]; 
    assign layer_0[2339] = ~(in[946] ^ in[931]); 
    assign layer_0[2340] = ~(in[925] | in[902]); 
    assign layer_0[2341] = ~(in[418] ^ in[486]); 
    assign layer_0[2342] = in[905] | in[598]; 
    assign layer_0[2343] = ~in[730]; 
    assign layer_0[2344] = in[36] ^ in[31]; 
    assign layer_0[2345] = in[520] ^ in[532]; 
    assign layer_0[2346] = in[339]; 
    assign layer_0[2347] = in[197] & ~in[126]; 
    assign layer_0[2348] = ~in[857] | (in[923] & in[857]); 
    assign layer_0[2349] = 1'b1; 
    assign layer_0[2350] = in[731] & in[439]; 
    assign layer_0[2351] = ~(in[904] | in[4]); 
    assign layer_0[2352] = ~(in[1003] ^ in[675]); 
    assign layer_0[2353] = in[431] ^ in[953]; 
    assign layer_0[2354] = ~(in[610] | in[529]); 
    assign layer_0[2355] = ~(in[499] ^ in[371]); 
    assign layer_0[2356] = ~(in[268] ^ in[235]); 
    assign layer_0[2357] = ~(in[921] ^ in[340]); 
    assign layer_0[2358] = ~(in[568] ^ in[796]); 
    assign layer_0[2359] = in[869]; 
    assign layer_0[2360] = in[968] ^ in[12]; 
    assign layer_0[2361] = in[702] & ~in[61]; 
    assign layer_0[2362] = in[908] ^ in[444]; 
    assign layer_0[2363] = in[290] & ~in[403]; 
    assign layer_0[2364] = in[759]; 
    assign layer_0[2365] = ~(in[395] & in[620]); 
    assign layer_0[2366] = ~(in[904] ^ in[935]); 
    assign layer_0[2367] = ~in[593]; 
    assign layer_0[2368] = in[175] ^ in[952]; 
    assign layer_0[2369] = ~(in[763] ^ in[156]); 
    assign layer_0[2370] = ~(in[629] ^ in[54]); 
    assign layer_0[2371] = ~in[359] | (in[553] & in[359]); 
    assign layer_0[2372] = ~(in[324] & in[512]); 
    assign layer_0[2373] = ~(in[843] | in[935]); 
    assign layer_0[2374] = ~in[740]; 
    assign layer_0[2375] = ~in[265] | (in[795] & in[265]); 
    assign layer_0[2376] = ~(in[239] & in[329]); 
    assign layer_0[2377] = in[493] ^ in[715]; 
    assign layer_0[2378] = ~(in[878] & in[669]); 
    assign layer_0[2379] = in[501]; 
    assign layer_0[2380] = ~(in[296] | in[722]); 
    assign layer_0[2381] = ~(in[1004] ^ in[632]); 
    assign layer_0[2382] = ~in[12]; 
    assign layer_0[2383] = 1'b0; 
    assign layer_0[2384] = in[388] & in[756]; 
    assign layer_0[2385] = ~in[569] | (in[779] & in[569]); 
    assign layer_0[2386] = ~(in[871] ^ in[872]); 
    assign layer_0[2387] = ~(in[350] ^ in[701]); 
    assign layer_0[2388] = ~(in[225] ^ in[508]); 
    assign layer_0[2389] = ~in[1013] | (in[573] & in[1013]); 
    assign layer_0[2390] = ~(in[67] & in[262]); 
    assign layer_0[2391] = in[771]; 
    assign layer_0[2392] = ~(in[364] ^ in[180]); 
    assign layer_0[2393] = in[915] ^ in[913]; 
    assign layer_0[2394] = ~in[83] | (in[905] & in[83]); 
    assign layer_0[2395] = ~(in[757] ^ in[740]); 
    assign layer_0[2396] = ~(in[995] ^ in[417]); 
    assign layer_0[2397] = ~(in[196] & in[377]); 
    assign layer_0[2398] = in[9] & ~in[791]; 
    assign layer_0[2399] = in[677] ^ in[635]; 
    assign layer_0[2400] = in[164] & ~in[702]; 
    assign layer_0[2401] = in[43] & in[665]; 
    assign layer_0[2402] = ~in[347]; 
    assign layer_0[2403] = in[190] & ~in[861]; 
    assign layer_0[2404] = in[841] & in[986]; 
    assign layer_0[2405] = in[583] ^ in[476]; 
    assign layer_0[2406] = in[319]; 
    assign layer_0[2407] = ~in[440]; 
    assign layer_0[2408] = in[824] & ~in[667]; 
    assign layer_0[2409] = ~in[872] | (in[541] & in[872]); 
    assign layer_0[2410] = ~(in[654] ^ in[741]); 
    assign layer_0[2411] = ~(in[769] ^ in[520]); 
    assign layer_0[2412] = in[855] & ~in[776]; 
    assign layer_0[2413] = ~(in[755] ^ in[599]); 
    assign layer_0[2414] = ~(in[260] ^ in[62]); 
    assign layer_0[2415] = 1'b1; 
    assign layer_0[2416] = ~(in[740] ^ in[965]); 
    assign layer_0[2417] = ~in[920]; 
    assign layer_0[2418] = ~(in[937] ^ in[450]); 
    assign layer_0[2419] = ~(in[260] & in[474]); 
    assign layer_0[2420] = ~in[143]; 
    assign layer_0[2421] = ~(in[857] ^ in[874]); 
    assign layer_0[2422] = in[969]; 
    assign layer_0[2423] = in[1000] ^ in[1001]; 
    assign layer_0[2424] = in[473] | in[843]; 
    assign layer_0[2425] = ~(in[981] ^ in[982]); 
    assign layer_0[2426] = ~(in[432] ^ in[21]); 
    assign layer_0[2427] = in[569]; 
    assign layer_0[2428] = ~(in[935] | in[887]); 
    assign layer_0[2429] = ~in[979] | (in[979] & in[589]); 
    assign layer_0[2430] = ~(in[313] ^ in[588]); 
    assign layer_0[2431] = ~(in[332] ^ in[449]); 
    assign layer_0[2432] = ~(in[968] ^ in[280]); 
    assign layer_0[2433] = ~in[742]; 
    assign layer_0[2434] = in[293] & in[83]; 
    assign layer_0[2435] = ~(in[254] | in[677]); 
    assign layer_0[2436] = in[227] ^ in[947]; 
    assign layer_0[2437] = in[842] ^ in[548]; 
    assign layer_0[2438] = ~(in[692] ^ in[519]); 
    assign layer_0[2439] = in[90] & in[178]; 
    assign layer_0[2440] = in[506] & ~in[95]; 
    assign layer_0[2441] = in[982]; 
    assign layer_0[2442] = ~(in[920] | in[722]); 
    assign layer_0[2443] = in[335] ^ in[711]; 
    assign layer_0[2444] = in[914] | in[811]; 
    assign layer_0[2445] = in[9] & in[151]; 
    assign layer_0[2446] = ~(in[588] ^ in[878]); 
    assign layer_0[2447] = ~(in[680] ^ in[632]); 
    assign layer_0[2448] = in[323] ^ in[708]; 
    assign layer_0[2449] = in[746] ^ in[5]; 
    assign layer_0[2450] = ~in[710]; 
    assign layer_0[2451] = ~in[851]; 
    assign layer_0[2452] = in[662] & ~in[899]; 
    assign layer_0[2453] = ~(in[511] ^ in[839]); 
    assign layer_0[2454] = ~in[596] | (in[583] & in[596]); 
    assign layer_0[2455] = ~in[101]; 
    assign layer_0[2456] = ~(in[666] ^ in[751]); 
    assign layer_0[2457] = ~in[141] | (in[141] & in[949]); 
    assign layer_0[2458] = ~in[98]; 
    assign layer_0[2459] = ~in[948] | (in[948] & in[872]); 
    assign layer_0[2460] = ~(in[628] ^ in[286]); 
    assign layer_0[2461] = ~in[583] | (in[583] & in[843]); 
    assign layer_0[2462] = in[966] & ~in[776]; 
    assign layer_0[2463] = ~(in[58] ^ in[397]); 
    assign layer_0[2464] = in[127] ^ in[13]; 
    assign layer_0[2465] = ~(in[477] ^ in[351]); 
    assign layer_0[2466] = ~(in[853] | in[815]); 
    assign layer_0[2467] = ~in[598]; 
    assign layer_0[2468] = ~(in[495] ^ in[861]); 
    assign layer_0[2469] = in[188] & ~in[916]; 
    assign layer_0[2470] = ~(in[551] ^ in[483]); 
    assign layer_0[2471] = in[873] ^ in[837]; 
    assign layer_0[2472] = ~in[316]; 
    assign layer_0[2473] = ~(in[227] ^ in[983]); 
    assign layer_0[2474] = ~(in[403] | in[571]); 
    assign layer_0[2475] = ~in[398] | (in[398] & in[729]); 
    assign layer_0[2476] = ~(in[14] ^ in[174]); 
    assign layer_0[2477] = ~in[602] | (in[602] & in[872]); 
    assign layer_0[2478] = in[387]; 
    assign layer_0[2479] = ~(in[1017] ^ in[920]); 
    assign layer_0[2480] = ~in[221] | (in[637] & in[221]); 
    assign layer_0[2481] = in[869] ^ in[870]; 
    assign layer_0[2482] = in[1002]; 
    assign layer_0[2483] = in[376] & in[477]; 
    assign layer_0[2484] = in[539]; 
    assign layer_0[2485] = ~(in[535] ^ in[923]); 
    assign layer_0[2486] = ~in[234]; 
    assign layer_0[2487] = ~in[518]; 
    assign layer_0[2488] = in[482] | in[338]; 
    assign layer_0[2489] = ~(in[168] ^ in[1018]); 
    assign layer_0[2490] = in[912] ^ in[934]; 
    assign layer_0[2491] = ~(in[519] ^ in[744]); 
    assign layer_0[2492] = ~(in[783] ^ in[707]); 
    assign layer_0[2493] = ~in[568]; 
    assign layer_0[2494] = ~in[55] | (in[55] & in[673]); 
    assign layer_0[2495] = ~in[938] | (in[719] & in[938]); 
    assign layer_0[2496] = in[110] & ~in[628]; 
    assign layer_0[2497] = in[1002] ^ in[274]; 
    assign layer_0[2498] = ~(in[457] ^ in[494]); 
    assign layer_0[2499] = in[286] ^ in[870]; 
    assign layer_0[2500] = ~(in[843] | in[867]); 
    assign layer_0[2501] = in[636] & ~in[737]; 
    assign layer_0[2502] = ~in[707] | (in[986] & in[707]); 
    assign layer_0[2503] = ~in[462]; 
    assign layer_0[2504] = ~in[904]; 
    assign layer_0[2505] = ~(in[719] ^ in[621]); 
    assign layer_0[2506] = ~(in[820] & in[216]); 
    assign layer_0[2507] = in[679] ^ in[312]; 
    assign layer_0[2508] = ~(in[931] ^ in[930]); 
    assign layer_0[2509] = ~in[18]; 
    assign layer_0[2510] = in[697] | in[626]; 
    assign layer_0[2511] = in[482] ^ in[761]; 
    assign layer_0[2512] = in[226] ^ in[28]; 
    assign layer_0[2513] = in[868] ^ in[580]; 
    assign layer_0[2514] = in[460] & ~in[126]; 
    assign layer_0[2515] = ~in[118] | (in[118] & in[753]); 
    assign layer_0[2516] = in[606] | in[552]; 
    assign layer_0[2517] = in[577]; 
    assign layer_0[2518] = ~(in[126] & in[68]); 
    assign layer_0[2519] = ~in[941]; 
    assign layer_0[2520] = ~in[593]; 
    assign layer_0[2521] = in[1015] & in[646]; 
    assign layer_0[2522] = ~(in[708] ^ in[243]); 
    assign layer_0[2523] = in[904]; 
    assign layer_0[2524] = in[482] ^ in[309]; 
    assign layer_0[2525] = in[298] ^ in[210]; 
    assign layer_0[2526] = in[838] ^ in[934]; 
    assign layer_0[2527] = in[845] ^ in[70]; 
    assign layer_0[2528] = ~(in[11] ^ in[884]); 
    assign layer_0[2529] = in[504] & ~in[609]; 
    assign layer_0[2530] = in[871] & in[983]; 
    assign layer_0[2531] = in[286] ^ in[399]; 
    assign layer_0[2532] = in[788] ^ in[696]; 
    assign layer_0[2533] = in[547] & ~in[698]; 
    assign layer_0[2534] = in[1018] | in[532]; 
    assign layer_0[2535] = in[946] ^ in[930]; 
    assign layer_0[2536] = ~in[963] | (in[963] & in[288]); 
    assign layer_0[2537] = in[688] ^ in[62]; 
    assign layer_0[2538] = ~in[71] | (in[71] & in[456]); 
    assign layer_0[2539] = ~(in[954] ^ in[533]); 
    assign layer_0[2540] = in[987] | in[262]; 
    assign layer_0[2541] = in[165] & in[216]; 
    assign layer_0[2542] = in[473] & in[938]; 
    assign layer_0[2543] = ~in[758] | (in[858] & in[758]); 
    assign layer_0[2544] = in[224]; 
    assign layer_0[2545] = in[662] ^ in[626]; 
    assign layer_0[2546] = in[660] | in[548]; 
    assign layer_0[2547] = in[937] ^ in[911]; 
    assign layer_0[2548] = ~(in[223] ^ in[131]); 
    assign layer_0[2549] = ~in[391] | (in[391] & in[459]); 
    assign layer_0[2550] = in[690] ^ in[307]; 
    assign layer_0[2551] = ~(in[826] ^ in[825]); 
    assign layer_0[2552] = in[581] & in[507]; 
    assign layer_0[2553] = in[837] ^ in[570]; 
    assign layer_0[2554] = in[976] & ~in[924]; 
    assign layer_0[2555] = in[869] & ~in[986]; 
    assign layer_0[2556] = ~(in[483] ^ in[950]); 
    assign layer_0[2557] = ~(in[371] ^ in[100]); 
    assign layer_0[2558] = ~in[850] | (in[850] & in[319]); 
    assign layer_0[2559] = in[520] ^ in[668]; 
    assign layer_0[2560] = in[840] ^ in[208]; 
    assign layer_0[2561] = in[357] & ~in[960]; 
    assign layer_0[2562] = in[930] | in[641]; 
    assign layer_0[2563] = ~(in[578] ^ in[614]); 
    assign layer_0[2564] = ~in[569]; 
    assign layer_0[2565] = in[220] & in[586]; 
    assign layer_0[2566] = ~in[982] | (in[844] & in[982]); 
    assign layer_0[2567] = ~(in[520] & in[823]); 
    assign layer_0[2568] = in[790]; 
    assign layer_0[2569] = in[397] & in[306]; 
    assign layer_0[2570] = ~in[931]; 
    assign layer_0[2571] = ~(in[162] ^ in[235]); 
    assign layer_0[2572] = in[73] & ~in[952]; 
    assign layer_0[2573] = in[479] | in[628]; 
    assign layer_0[2574] = in[66] ^ in[451]; 
    assign layer_0[2575] = ~in[20] | (in[20] & in[130]); 
    assign layer_0[2576] = ~in[51]; 
    assign layer_0[2577] = ~(in[317] ^ in[652]); 
    assign layer_0[2578] = in[484] | in[822]; 
    assign layer_0[2579] = in[509] ^ in[966]; 
    assign layer_0[2580] = ~(in[301] ^ in[447]); 
    assign layer_0[2581] = ~(in[398] ^ in[959]); 
    assign layer_0[2582] = ~in[719]; 
    assign layer_0[2583] = in[931] ^ in[498]; 
    assign layer_0[2584] = in[44] | in[331]; 
    assign layer_0[2585] = in[429]; 
    assign layer_0[2586] = in[936] & ~in[709]; 
    assign layer_0[2587] = ~in[519]; 
    assign layer_0[2588] = ~in[776] | (in[315] & in[776]); 
    assign layer_0[2589] = ~(in[790] ^ in[809]); 
    assign layer_0[2590] = ~in[610] | (in[610] & in[10]); 
    assign layer_0[2591] = ~in[67] | (in[574] & in[67]); 
    assign layer_0[2592] = ~in[616] | (in[616] & in[341]); 
    assign layer_0[2593] = in[858]; 
    assign layer_0[2594] = ~(in[615] & in[465]); 
    assign layer_0[2595] = in[433]; 
    assign layer_0[2596] = in[520]; 
    assign layer_0[2597] = ~(in[1019] ^ in[874]); 
    assign layer_0[2598] = ~in[309]; 
    assign layer_0[2599] = in[821] ^ in[704]; 
    assign layer_0[2600] = in[822] ^ in[776]; 
    assign layer_0[2601] = ~in[429] | (in[429] & in[481]); 
    assign layer_0[2602] = ~(in[360] & in[788]); 
    assign layer_0[2603] = ~in[587] | (in[587] & in[241]); 
    assign layer_0[2604] = ~(in[897] | in[582]); 
    assign layer_0[2605] = ~(in[289] | in[483]); 
    assign layer_0[2606] = ~(in[997] ^ in[931]); 
    assign layer_0[2607] = in[792] ^ in[579]; 
    assign layer_0[2608] = ~(in[844] | in[241]); 
    assign layer_0[2609] = ~(in[688] | in[268]); 
    assign layer_0[2610] = in[476] ^ in[1003]; 
    assign layer_0[2611] = in[852] | in[936]; 
    assign layer_0[2612] = ~(in[877] | in[77]); 
    assign layer_0[2613] = ~(in[694] ^ in[388]); 
    assign layer_0[2614] = ~in[261] | (in[261] & in[264]); 
    assign layer_0[2615] = in[889] | in[627]; 
    assign layer_0[2616] = in[865]; 
    assign layer_0[2617] = ~(in[928] ^ in[892]); 
    assign layer_0[2618] = ~(in[692] ^ in[19]); 
    assign layer_0[2619] = ~in[536] | (in[872] & in[536]); 
    assign layer_0[2620] = ~in[603] | (in[333] & in[603]); 
    assign layer_0[2621] = ~(in[266] & in[345]); 
    assign layer_0[2622] = in[524] | in[435]; 
    assign layer_0[2623] = in[565] ^ in[276]; 
    assign layer_0[2624] = in[835] & ~in[243]; 
    assign layer_0[2625] = in[619] ^ in[178]; 
    assign layer_0[2626] = ~(in[277] ^ in[382]); 
    assign layer_0[2627] = in[483] ^ in[109]; 
    assign layer_0[2628] = ~in[502] | (in[502] & in[510]); 
    assign layer_0[2629] = ~(in[616] ^ in[622]); 
    assign layer_0[2630] = ~(in[569] & in[250]); 
    assign layer_0[2631] = in[149]; 
    assign layer_0[2632] = ~in[659] | (in[659] & in[134]); 
    assign layer_0[2633] = in[441] & ~in[35]; 
    assign layer_0[2634] = ~in[449]; 
    assign layer_0[2635] = in[732]; 
    assign layer_0[2636] = ~(in[429] & in[125]); 
    assign layer_0[2637] = in[279]; 
    assign layer_0[2638] = ~(in[532] | in[382]); 
    assign layer_0[2639] = ~in[647] | (in[647] & in[836]); 
    assign layer_0[2640] = ~in[193] | (in[325] & in[193]); 
    assign layer_0[2641] = in[145]; 
    assign layer_0[2642] = ~in[944]; 
    assign layer_0[2643] = in[936]; 
    assign layer_0[2644] = ~(in[730] ^ in[954]); 
    assign layer_0[2645] = ~(in[890] ^ in[459]); 
    assign layer_0[2646] = ~(in[18] ^ in[519]); 
    assign layer_0[2647] = in[302] & ~in[354]; 
    assign layer_0[2648] = in[5]; 
    assign layer_0[2649] = ~(in[823] ^ in[82]); 
    assign layer_0[2650] = ~in[210]; 
    assign layer_0[2651] = ~(in[921] ^ in[985]); 
    assign layer_0[2652] = in[706] ^ in[862]; 
    assign layer_0[2653] = ~(in[159] | in[964]); 
    assign layer_0[2654] = ~(in[950] & in[152]); 
    assign layer_0[2655] = in[116] ^ in[393]; 
    assign layer_0[2656] = ~(in[3] ^ in[429]); 
    assign layer_0[2657] = in[905]; 
    assign layer_0[2658] = in[410] & in[759]; 
    assign layer_0[2659] = ~in[581] | (in[581] & in[747]); 
    assign layer_0[2660] = in[982] ^ in[597]; 
    assign layer_0[2661] = in[205] & in[856]; 
    assign layer_0[2662] = ~in[317] | (in[317] & in[3]); 
    assign layer_0[2663] = ~in[859] | (in[859] & in[917]); 
    assign layer_0[2664] = ~(in[432] ^ in[253]); 
    assign layer_0[2665] = in[885] ^ in[658]; 
    assign layer_0[2666] = ~in[907]; 
    assign layer_0[2667] = in[386] ^ in[266]; 
    assign layer_0[2668] = in[731] | in[794]; 
    assign layer_0[2669] = ~(in[657] | in[627]); 
    assign layer_0[2670] = in[461] & in[443]; 
    assign layer_0[2671] = ~in[899]; 
    assign layer_0[2672] = in[638] & in[651]; 
    assign layer_0[2673] = ~(in[825] ^ in[842]); 
    assign layer_0[2674] = ~in[321] | (in[321] & in[963]); 
    assign layer_0[2675] = in[904] | in[776]; 
    assign layer_0[2676] = in[322] ^ in[658]; 
    assign layer_0[2677] = ~(in[809] ^ in[808]); 
    assign layer_0[2678] = ~in[373] | (in[373] & in[364]); 
    assign layer_0[2679] = ~in[1010] | (in[190] & in[1010]); 
    assign layer_0[2680] = ~(in[254] ^ in[571]); 
    assign layer_0[2681] = in[421] | in[181]; 
    assign layer_0[2682] = in[1022] ^ in[858]; 
    assign layer_0[2683] = ~(in[908] & in[188]); 
    assign layer_0[2684] = in[387] ^ in[572]; 
    assign layer_0[2685] = in[959] | in[904]; 
    assign layer_0[2686] = ~(in[823] ^ in[889]); 
    assign layer_0[2687] = ~in[890]; 
    assign layer_0[2688] = in[266]; 
    assign layer_0[2689] = ~(in[895] | in[278]); 
    assign layer_0[2690] = in[626] ^ in[253]; 
    assign layer_0[2691] = in[368] ^ in[685]; 
    assign layer_0[2692] = in[813] | in[1005]; 
    assign layer_0[2693] = 1'b0; 
    assign layer_0[2694] = in[819] & ~in[398]; 
    assign layer_0[2695] = in[321] & in[808]; 
    assign layer_0[2696] = ~in[307] | (in[307] & in[193]); 
    assign layer_0[2697] = ~(in[539] & in[469]); 
    assign layer_0[2698] = ~in[259] | (in[188] & in[259]); 
    assign layer_0[2699] = in[734] & ~in[86]; 
    assign layer_0[2700] = ~(in[241] ^ in[312]); 
    assign layer_0[2701] = ~in[26]; 
    assign layer_0[2702] = in[226]; 
    assign layer_0[2703] = ~(in[923] ^ in[844]); 
    assign layer_0[2704] = in[927] ^ in[623]; 
    assign layer_0[2705] = ~(in[161] ^ in[114]); 
    assign layer_0[2706] = ~(in[101] | in[986]); 
    assign layer_0[2707] = in[627] ^ in[931]; 
    assign layer_0[2708] = ~in[775]; 
    assign layer_0[2709] = in[241] ^ in[282]; 
    assign layer_0[2710] = ~in[516] | (in[516] & in[765]); 
    assign layer_0[2711] = ~(in[283] ^ in[181]); 
    assign layer_0[2712] = ~(in[250] | in[658]); 
    assign layer_0[2713] = in[650] ^ in[754]; 
    assign layer_0[2714] = ~in[690] | (in[38] & in[690]); 
    assign layer_0[2715] = in[5] & ~in[459]; 
    assign layer_0[2716] = in[883] & in[876]; 
    assign layer_0[2717] = in[314] & ~in[378]; 
    assign layer_0[2718] = in[139] | in[432]; 
    assign layer_0[2719] = ~(in[589] ^ in[741]); 
    assign layer_0[2720] = ~(in[61] ^ in[315]); 
    assign layer_0[2721] = ~in[930] | (in[930] & in[977]); 
    assign layer_0[2722] = ~(in[440] & in[997]); 
    assign layer_0[2723] = in[940] & in[174]; 
    assign layer_0[2724] = ~(in[551] & in[263]); 
    assign layer_0[2725] = in[572] ^ in[605]; 
    assign layer_0[2726] = in[236] ^ in[857]; 
    assign layer_0[2727] = ~in[19] | (in[19] & in[434]); 
    assign layer_0[2728] = in[238] ^ in[792]; 
    assign layer_0[2729] = in[467]; 
    assign layer_0[2730] = in[890]; 
    assign layer_0[2731] = ~(in[505] & in[356]); 
    assign layer_0[2732] = ~(in[799] ^ in[732]); 
    assign layer_0[2733] = in[155] & ~in[250]; 
    assign layer_0[2734] = in[365] ^ in[13]; 
    assign layer_0[2735] = ~in[19] | (in[19] & in[919]); 
    assign layer_0[2736] = ~in[391]; 
    assign layer_0[2737] = in[323] & in[725]; 
    assign layer_0[2738] = ~in[598] | (in[598] & in[924]); 
    assign layer_0[2739] = ~(in[574] | in[479]); 
    assign layer_0[2740] = in[614] & ~in[337]; 
    assign layer_0[2741] = in[632] & ~in[38]; 
    assign layer_0[2742] = ~(in[937] ^ in[648]); 
    assign layer_0[2743] = in[499] & in[607]; 
    assign layer_0[2744] = ~(in[552] & in[260]); 
    assign layer_0[2745] = in[571] ^ in[130]; 
    assign layer_0[2746] = in[413] ^ in[13]; 
    assign layer_0[2747] = ~(in[299] & in[605]); 
    assign layer_0[2748] = ~in[172] | (in[927] & in[172]); 
    assign layer_0[2749] = ~(in[381] & in[317]); 
    assign layer_0[2750] = in[611] | in[239]; 
    assign layer_0[2751] = in[762] ^ in[774]; 
    assign layer_0[2752] = in[536] ^ in[680]; 
    assign layer_0[2753] = ~(in[1008] | in[920]); 
    assign layer_0[2754] = ~in[894] | (in[742] & in[894]); 
    assign layer_0[2755] = ~(in[788] ^ in[178]); 
    assign layer_0[2756] = ~in[156] | (in[156] & in[95]); 
    assign layer_0[2757] = ~(in[1000] ^ in[612]); 
    assign layer_0[2758] = ~(in[122] & in[585]); 
    assign layer_0[2759] = in[987] ^ in[873]; 
    assign layer_0[2760] = in[578] & ~in[515]; 
    assign layer_0[2761] = in[763]; 
    assign layer_0[2762] = ~(in[59] | in[526]); 
    assign layer_0[2763] = in[65] | in[838]; 
    assign layer_0[2764] = in[952]; 
    assign layer_0[2765] = ~(in[637] ^ in[954]); 
    assign layer_0[2766] = 1'b0; 
    assign layer_0[2767] = ~(in[256] | in[951]); 
    assign layer_0[2768] = in[922] | in[143]; 
    assign layer_0[2769] = ~(in[883] | in[553]); 
    assign layer_0[2770] = in[409] & ~in[263]; 
    assign layer_0[2771] = ~in[51] | (in[51] & in[30]); 
    assign layer_0[2772] = in[870]; 
    assign layer_0[2773] = ~in[936]; 
    assign layer_0[2774] = in[598] & ~in[829]; 
    assign layer_0[2775] = ~(in[766] | in[94]); 
    assign layer_0[2776] = ~(in[706] ^ in[988]); 
    assign layer_0[2777] = ~(in[974] ^ in[662]); 
    assign layer_0[2778] = ~(in[287] | in[566]); 
    assign layer_0[2779] = ~in[593] | (in[984] & in[593]); 
    assign layer_0[2780] = in[501] & ~in[558]; 
    assign layer_0[2781] = in[618] & ~in[748]; 
    assign layer_0[2782] = in[812] ^ in[828]; 
    assign layer_0[2783] = ~in[340]; 
    assign layer_0[2784] = in[565] ^ in[555]; 
    assign layer_0[2785] = ~in[955] | (in[623] & in[955]); 
    assign layer_0[2786] = ~(in[935] ^ in[50]); 
    assign layer_0[2787] = in[91] ^ in[670]; 
    assign layer_0[2788] = ~in[618] | (in[389] & in[618]); 
    assign layer_0[2789] = ~in[757] | (in[757] & in[605]); 
    assign layer_0[2790] = in[646] & ~in[249]; 
    assign layer_0[2791] = in[135] ^ in[449]; 
    assign layer_0[2792] = in[635]; 
    assign layer_0[2793] = in[596] ^ in[661]; 
    assign layer_0[2794] = in[396] & in[399]; 
    assign layer_0[2795] = in[365] | in[334]; 
    assign layer_0[2796] = ~(in[1018] ^ in[844]); 
    assign layer_0[2797] = ~(in[603] | in[538]); 
    assign layer_0[2798] = ~in[632] | (in[224] & in[632]); 
    assign layer_0[2799] = ~(in[970] ^ in[444]); 
    assign layer_0[2800] = in[587] ^ in[326]; 
    assign layer_0[2801] = ~(in[966] ^ in[967]); 
    assign layer_0[2802] = ~(in[628] | in[96]); 
    assign layer_0[2803] = in[664] & ~in[531]; 
    assign layer_0[2804] = ~in[157] | (in[157] & in[499]); 
    assign layer_0[2805] = ~(in[859] | in[211]); 
    assign layer_0[2806] = ~(in[572] & in[551]); 
    assign layer_0[2807] = ~in[983] | (in[966] & in[983]); 
    assign layer_0[2808] = in[203] & ~in[755]; 
    assign layer_0[2809] = in[605] ^ in[570]; 
    assign layer_0[2810] = ~(in[624] | in[853]); 
    assign layer_0[2811] = in[718] ^ in[729]; 
    assign layer_0[2812] = in[902] | in[904]; 
    assign layer_0[2813] = in[824] & ~in[800]; 
    assign layer_0[2814] = in[46] | in[1016]; 
    assign layer_0[2815] = in[846] & ~in[547]; 
    assign layer_0[2816] = in[146] & ~in[21]; 
    assign layer_0[2817] = ~(in[194] ^ in[394]); 
    assign layer_0[2818] = in[445] ^ in[747]; 
    assign layer_0[2819] = ~in[277] | (in[277] & in[765]); 
    assign layer_0[2820] = in[578] | in[480]; 
    assign layer_0[2821] = in[1005] ^ in[698]; 
    assign layer_0[2822] = ~(in[413] | in[523]); 
    assign layer_0[2823] = in[968] | in[698]; 
    assign layer_0[2824] = ~(in[535] ^ in[569]); 
    assign layer_0[2825] = ~in[322] | (in[450] & in[322]); 
    assign layer_0[2826] = ~in[951]; 
    assign layer_0[2827] = ~in[934] | (in[759] & in[934]); 
    assign layer_0[2828] = in[143] ^ in[9]; 
    assign layer_0[2829] = ~in[1009] | (in[531] & in[1009]); 
    assign layer_0[2830] = in[600] & ~in[629]; 
    assign layer_0[2831] = ~(in[373] ^ in[450]); 
    assign layer_0[2832] = in[457] & in[830]; 
    assign layer_0[2833] = in[939] & ~in[737]; 
    assign layer_0[2834] = ~(in[685] ^ in[583]); 
    assign layer_0[2835] = in[784]; 
    assign layer_0[2836] = in[431]; 
    assign layer_0[2837] = ~in[526]; 
    assign layer_0[2838] = ~(in[390] ^ in[716]); 
    assign layer_0[2839] = ~(in[950] ^ in[242]); 
    assign layer_0[2840] = 1'b0; 
    assign layer_0[2841] = in[855] ^ in[312]; 
    assign layer_0[2842] = in[869] ^ in[858]; 
    assign layer_0[2843] = in[646] & ~in[14]; 
    assign layer_0[2844] = in[714] & ~in[533]; 
    assign layer_0[2845] = ~(in[914] ^ in[483]); 
    assign layer_0[2846] = ~in[169]; 
    assign layer_0[2847] = in[54] & ~in[33]; 
    assign layer_0[2848] = in[663]; 
    assign layer_0[2849] = ~(in[918] ^ in[987]); 
    assign layer_0[2850] = in[691] ^ in[195]; 
    assign layer_0[2851] = ~(in[339] | in[644]); 
    assign layer_0[2852] = ~(in[2] | in[354]); 
    assign layer_0[2853] = ~(in[939] ^ in[909]); 
    assign layer_0[2854] = ~in[234]; 
    assign layer_0[2855] = ~(in[624] | in[209]); 
    assign layer_0[2856] = ~in[730]; 
    assign layer_0[2857] = ~in[804]; 
    assign layer_0[2858] = in[139] & in[419]; 
    assign layer_0[2859] = ~in[266] | (in[266] & in[718]); 
    assign layer_0[2860] = ~(in[218] | in[680]); 
    assign layer_0[2861] = in[604]; 
    assign layer_0[2862] = in[870] ^ in[917]; 
    assign layer_0[2863] = in[930] & ~in[222]; 
    assign layer_0[2864] = in[710]; 
    assign layer_0[2865] = ~(in[141] | in[366]); 
    assign layer_0[2866] = ~(in[284] | in[950]); 
    assign layer_0[2867] = in[37]; 
    assign layer_0[2868] = in[57] ^ in[758]; 
    assign layer_0[2869] = in[781] & in[828]; 
    assign layer_0[2870] = ~(in[708] ^ in[509]); 
    assign layer_0[2871] = ~in[228] | (in[403] & in[228]); 
    assign layer_0[2872] = in[748]; 
    assign layer_0[2873] = ~(in[431] & in[945]); 
    assign layer_0[2874] = ~in[537] | (in[860] & in[537]); 
    assign layer_0[2875] = in[222]; 
    assign layer_0[2876] = in[251] & ~in[988]; 
    assign layer_0[2877] = ~(in[287] | in[981]); 
    assign layer_0[2878] = ~in[878] | (in[878] & in[138]); 
    assign layer_0[2879] = in[517] & in[154]; 
    assign layer_0[2880] = in[156] | in[236]; 
    assign layer_0[2881] = in[549] & in[837]; 
    assign layer_0[2882] = in[369] ^ in[874]; 
    assign layer_0[2883] = in[934]; 
    assign layer_0[2884] = in[972] & in[265]; 
    assign layer_0[2885] = in[520] & ~in[732]; 
    assign layer_0[2886] = ~(in[933] ^ in[30]); 
    assign layer_0[2887] = in[683] ^ in[590]; 
    assign layer_0[2888] = ~in[884]; 
    assign layer_0[2889] = in[160] ^ in[885]; 
    assign layer_0[2890] = ~in[252] | (in[155] & in[252]); 
    assign layer_0[2891] = ~in[901] | (in[367] & in[901]); 
    assign layer_0[2892] = ~in[252]; 
    assign layer_0[2893] = ~in[308]; 
    assign layer_0[2894] = ~(in[597] ^ in[418]); 
    assign layer_0[2895] = ~(in[476] ^ in[644]); 
    assign layer_0[2896] = in[702] ^ in[165]; 
    assign layer_0[2897] = in[427] & ~in[894]; 
    assign layer_0[2898] = in[701] & ~in[230]; 
    assign layer_0[2899] = in[1004]; 
    assign layer_0[2900] = in[693]; 
    assign layer_0[2901] = in[364] ^ in[436]; 
    assign layer_0[2902] = ~(in[284] ^ in[792]); 
    assign layer_0[2903] = ~in[265] | (in[28] & in[265]); 
    assign layer_0[2904] = ~in[456] | (in[1001] & in[456]); 
    assign layer_0[2905] = ~in[319]; 
    assign layer_0[2906] = in[351] ^ in[451]; 
    assign layer_0[2907] = ~in[747] | (in[642] & in[747]); 
    assign layer_0[2908] = in[963] & ~in[209]; 
    assign layer_0[2909] = ~in[792]; 
    assign layer_0[2910] = ~(in[595] | in[792]); 
    assign layer_0[2911] = ~(in[659] ^ in[227]); 
    assign layer_0[2912] = in[459] & in[485]; 
    assign layer_0[2913] = 1'b1; 
    assign layer_0[2914] = ~in[985]; 
    assign layer_0[2915] = 1'b0; 
    assign layer_0[2916] = in[932] & ~in[672]; 
    assign layer_0[2917] = ~(in[651] & in[229]); 
    assign layer_0[2918] = ~in[295] | (in[295] & in[282]); 
    assign layer_0[2919] = in[629] ^ in[251]; 
    assign layer_0[2920] = in[687] & ~in[38]; 
    assign layer_0[2921] = ~(in[252] ^ in[958]); 
    assign layer_0[2922] = ~in[103] | (in[999] & in[103]); 
    assign layer_0[2923] = in[441] & ~in[328]; 
    assign layer_0[2924] = in[618] ^ in[658]; 
    assign layer_0[2925] = ~(in[999] | in[667]); 
    assign layer_0[2926] = ~(in[11] ^ in[193]); 
    assign layer_0[2927] = in[910] ^ in[688]; 
    assign layer_0[2928] = in[92] ^ in[640]; 
    assign layer_0[2929] = in[743] | in[973]; 
    assign layer_0[2930] = ~(in[508] ^ in[920]); 
    assign layer_0[2931] = in[638] & ~in[680]; 
    assign layer_0[2932] = 1'b0; 
    assign layer_0[2933] = in[627]; 
    assign layer_0[2934] = in[739] ^ in[464]; 
    assign layer_0[2935] = in[759] ^ in[519]; 
    assign layer_0[2936] = ~(in[821] ^ in[266]); 
    assign layer_0[2937] = in[865] | in[86]; 
    assign layer_0[2938] = in[482] ^ in[853]; 
    assign layer_0[2939] = ~(in[326] ^ in[764]); 
    assign layer_0[2940] = ~in[702] | (in[319] & in[702]); 
    assign layer_0[2941] = in[738] & ~in[1002]; 
    assign layer_0[2942] = ~in[436] | (in[436] & in[604]); 
    assign layer_0[2943] = in[585] ^ in[757]; 
    assign layer_0[2944] = ~(in[459] & in[654]); 
    assign layer_0[2945] = in[358] | in[206]; 
    assign layer_0[2946] = ~in[912]; 
    assign layer_0[2947] = in[746] | in[617]; 
    assign layer_0[2948] = in[571]; 
    assign layer_0[2949] = in[499] ^ in[56]; 
    assign layer_0[2950] = in[537] & ~in[79]; 
    assign layer_0[2951] = ~(in[20] ^ in[947]); 
    assign layer_0[2952] = ~in[644] | (in[740] & in[644]); 
    assign layer_0[2953] = ~(in[869] ^ in[520]); 
    assign layer_0[2954] = ~in[180] | (in[180] & in[348]); 
    assign layer_0[2955] = ~in[363]; 
    assign layer_0[2956] = in[210] & ~in[286]; 
    assign layer_0[2957] = ~in[551] | (in[841] & in[551]); 
    assign layer_0[2958] = ~in[937]; 
    assign layer_0[2959] = ~(in[868] | in[575]); 
    assign layer_0[2960] = ~(in[757] ^ in[617]); 
    assign layer_0[2961] = in[246] & ~in[498]; 
    assign layer_0[2962] = ~(in[81] | in[533]); 
    assign layer_0[2963] = in[843] ^ in[703]; 
    assign layer_0[2964] = ~in[436] | (in[876] & in[436]); 
    assign layer_0[2965] = in[1008] | in[1010]; 
    assign layer_0[2966] = in[142] & ~in[289]; 
    assign layer_0[2967] = ~(in[346] ^ in[597]); 
    assign layer_0[2968] = in[396] ^ in[538]; 
    assign layer_0[2969] = ~in[1014] | (in[1014] & in[676]); 
    assign layer_0[2970] = ~(in[385] | in[84]); 
    assign layer_0[2971] = ~in[796] | (in[623] & in[796]); 
    assign layer_0[2972] = in[174] ^ in[694]; 
    assign layer_0[2973] = in[434] & in[836]; 
    assign layer_0[2974] = ~in[956]; 
    assign layer_0[2975] = ~in[633] | (in[633] & in[835]); 
    assign layer_0[2976] = ~(in[724] ^ in[595]); 
    assign layer_0[2977] = in[4] ^ in[131]; 
    assign layer_0[2978] = in[940]; 
    assign layer_0[2979] = ~(in[274] ^ in[934]); 
    assign layer_0[2980] = ~(in[1022] | in[277]); 
    assign layer_0[2981] = ~in[682] | (in[68] & in[682]); 
    assign layer_0[2982] = ~(in[652] ^ in[899]); 
    assign layer_0[2983] = in[867] ^ in[508]; 
    assign layer_0[2984] = in[716] ^ in[503]; 
    assign layer_0[2985] = in[306]; 
    assign layer_0[2986] = ~in[260] | (in[260] & in[908]); 
    assign layer_0[2987] = ~(in[595] & in[291]); 
    assign layer_0[2988] = in[875] ^ in[318]; 
    assign layer_0[2989] = ~in[672] | (in[672] & in[232]); 
    assign layer_0[2990] = ~(in[595] | in[971]); 
    assign layer_0[2991] = ~(in[124] ^ in[300]); 
    assign layer_0[2992] = in[819] | in[285]; 
    assign layer_0[2993] = in[500] ^ in[260]; 
    assign layer_0[2994] = ~in[190] | (in[190] & in[144]); 
    assign layer_0[2995] = in[952] & ~in[800]; 
    assign layer_0[2996] = ~(in[546] | in[598]); 
    assign layer_0[2997] = ~in[561]; 
    assign layer_0[2998] = ~(in[769] ^ in[201]); 
    assign layer_0[2999] = in[516]; 
    assign layer_0[3000] = ~in[915] | (in[507] & in[915]); 
    assign layer_0[3001] = ~in[263]; 
    assign layer_0[3002] = in[438] & ~in[755]; 
    assign layer_0[3003] = in[821] | in[68]; 
    assign layer_0[3004] = ~(in[926] ^ in[435]); 
    assign layer_0[3005] = ~in[296]; 
    assign layer_0[3006] = in[856] ^ in[602]; 
    assign layer_0[3007] = in[259] | in[826]; 
    assign layer_0[3008] = in[633] | in[906]; 
    assign layer_0[3009] = in[163] & ~in[1014]; 
    assign layer_0[3010] = 1'b0; 
    assign layer_0[3011] = in[932] ^ in[237]; 
    assign layer_0[3012] = ~(in[381] ^ in[29]); 
    assign layer_0[3013] = in[1017] ^ in[1016]; 
    assign layer_0[3014] = in[664] & ~in[34]; 
    assign layer_0[3015] = ~in[37] | (in[37] & in[624]); 
    assign layer_0[3016] = ~in[518] | (in[824] & in[518]); 
    assign layer_0[3017] = in[19]; 
    assign layer_0[3018] = in[956]; 
    assign layer_0[3019] = ~(in[11] ^ in[776]); 
    assign layer_0[3020] = in[641] & in[376]; 
    assign layer_0[3021] = ~in[613] | (in[613] & in[888]); 
    assign layer_0[3022] = ~(in[581] & in[548]); 
    assign layer_0[3023] = in[3]; 
    assign layer_0[3024] = ~in[78] | (in[78] & in[706]); 
    assign layer_0[3025] = in[694] ^ in[611]; 
    assign layer_0[3026] = in[284] ^ in[888]; 
    assign layer_0[3027] = ~(in[584] | in[282]); 
    assign layer_0[3028] = ~in[891] | (in[891] & in[267]); 
    assign layer_0[3029] = in[15] ^ in[594]; 
    assign layer_0[3030] = ~(in[348] ^ in[483]); 
    assign layer_0[3031] = ~in[941]; 
    assign layer_0[3032] = in[27]; 
    assign layer_0[3033] = ~(in[354] ^ in[353]); 
    assign layer_0[3034] = in[346] & ~in[511]; 
    assign layer_0[3035] = ~(in[333] ^ in[264]); 
    assign layer_0[3036] = in[691] | in[684]; 
    assign layer_0[3037] = ~(in[894] ^ in[21]); 
    assign layer_0[3038] = ~(in[677] & in[757]); 
    assign layer_0[3039] = ~(in[683] | in[272]); 
    assign layer_0[3040] = ~in[264] | (in[264] & in[207]); 
    assign layer_0[3041] = ~in[106] | (in[572] & in[106]); 
    assign layer_0[3042] = in[902] & ~in[221]; 
    assign layer_0[3043] = ~(in[253] ^ in[551]); 
    assign layer_0[3044] = ~in[163] | (in[163] & in[491]); 
    assign layer_0[3045] = in[709] & ~in[994]; 
    assign layer_0[3046] = ~(in[726] ^ in[804]); 
    assign layer_0[3047] = ~in[44] | (in[243] & in[44]); 
    assign layer_0[3048] = in[537] | in[545]; 
    assign layer_0[3049] = ~(in[614] ^ in[142]); 
    assign layer_0[3050] = ~(in[709] ^ in[465]); 
    assign layer_0[3051] = in[339] | in[348]; 
    assign layer_0[3052] = in[922] & ~in[554]; 
    assign layer_0[3053] = in[953] ^ in[473]; 
    assign layer_0[3054] = in[699]; 
    assign layer_0[3055] = ~in[836]; 
    assign layer_0[3056] = ~(in[968] ^ in[602]); 
    assign layer_0[3057] = ~in[638] | (in[638] & in[574]); 
    assign layer_0[3058] = in[62] ^ in[731]; 
    assign layer_0[3059] = in[572] ^ in[568]; 
    assign layer_0[3060] = in[402] | in[1014]; 
    assign layer_0[3061] = ~in[95]; 
    assign layer_0[3062] = in[179] ^ in[483]; 
    assign layer_0[3063] = in[166] | in[394]; 
    assign layer_0[3064] = in[104] & ~in[939]; 
    assign layer_0[3065] = ~in[652] | (in[652] & in[225]); 
    assign layer_0[3066] = in[759] ^ in[792]; 
    assign layer_0[3067] = ~in[47]; 
    assign layer_0[3068] = ~(in[464] & in[85]); 
    assign layer_0[3069] = in[101] & in[903]; 
    assign layer_0[3070] = in[217] ^ in[423]; 
    assign layer_0[3071] = in[976]; 
    assign layer_0[3072] = ~in[807]; 
    assign layer_0[3073] = ~in[579]; 
    assign layer_0[3074] = in[505] | in[904]; 
    assign layer_0[3075] = ~(in[8] | in[657]); 
    assign layer_0[3076] = ~in[90]; 
    assign layer_0[3077] = in[342] & ~in[886]; 
    assign layer_0[3078] = in[460] & ~in[31]; 
    assign layer_0[3079] = ~(in[600] ^ in[601]); 
    assign layer_0[3080] = ~in[920]; 
    assign layer_0[3081] = in[599] ^ in[983]; 
    assign layer_0[3082] = in[461] & ~in[847]; 
    assign layer_0[3083] = ~(in[600] ^ in[466]); 
    assign layer_0[3084] = in[869] ^ in[842]; 
    assign layer_0[3085] = ~in[963] | (in[564] & in[963]); 
    assign layer_0[3086] = in[857]; 
    assign layer_0[3087] = ~(in[507] ^ in[792]); 
    assign layer_0[3088] = in[729] ^ in[722]; 
    assign layer_0[3089] = in[686] & ~in[502]; 
    assign layer_0[3090] = in[520] & ~in[482]; 
    assign layer_0[3091] = ~in[476] | (in[476] & in[131]); 
    assign layer_0[3092] = in[992] | in[35]; 
    assign layer_0[3093] = ~in[593]; 
    assign layer_0[3094] = ~(in[935] ^ in[1018]); 
    assign layer_0[3095] = in[569] ^ in[568]; 
    assign layer_0[3096] = in[305] & in[1022]; 
    assign layer_0[3097] = ~in[252] | (in[364] & in[252]); 
    assign layer_0[3098] = ~in[730]; 
    assign layer_0[3099] = in[504] & ~in[952]; 
    assign layer_0[3100] = in[45] | in[581]; 
    assign layer_0[3101] = in[716] ^ in[473]; 
    assign layer_0[3102] = in[0] ^ in[681]; 
    assign layer_0[3103] = ~(in[308] ^ in[62]); 
    assign layer_0[3104] = in[76] ^ in[932]; 
    assign layer_0[3105] = ~(in[999] ^ in[922]); 
    assign layer_0[3106] = in[129]; 
    assign layer_0[3107] = in[960] ^ in[781]; 
    assign layer_0[3108] = in[823]; 
    assign layer_0[3109] = ~(in[878] ^ in[717]); 
    assign layer_0[3110] = in[375]; 
    assign layer_0[3111] = in[283] | in[815]; 
    assign layer_0[3112] = ~in[170] | (in[916] & in[170]); 
    assign layer_0[3113] = in[643]; 
    assign layer_0[3114] = ~(in[391] ^ in[934]); 
    assign layer_0[3115] = ~in[375]; 
    assign layer_0[3116] = in[777]; 
    assign layer_0[3117] = ~(in[760] ^ in[501]); 
    assign layer_0[3118] = ~in[42] | (in[553] & in[42]); 
    assign layer_0[3119] = in[853] & ~in[807]; 
    assign layer_0[3120] = in[861] ^ in[925]; 
    assign layer_0[3121] = ~(in[996] ^ in[632]); 
    assign layer_0[3122] = ~(in[732] ^ in[84]); 
    assign layer_0[3123] = in[730]; 
    assign layer_0[3124] = ~in[369] | (in[369] & in[66]); 
    assign layer_0[3125] = ~(in[276] ^ in[413]); 
    assign layer_0[3126] = in[604] ^ in[250]; 
    assign layer_0[3127] = in[191] & in[870]; 
    assign layer_0[3128] = in[114] ^ in[62]; 
    assign layer_0[3129] = ~(in[614] ^ in[955]); 
    assign layer_0[3130] = in[604] ^ in[348]; 
    assign layer_0[3131] = ~(in[24] ^ in[843]); 
    assign layer_0[3132] = ~in[504] | (in[504] & in[334]); 
    assign layer_0[3133] = in[839] ^ in[872]; 
    assign layer_0[3134] = in[7] ^ in[354]; 
    assign layer_0[3135] = ~in[708] | (in[545] & in[708]); 
    assign layer_0[3136] = in[842] ^ in[790]; 
    assign layer_0[3137] = in[679] & ~in[888]; 
    assign layer_0[3138] = in[262] & ~in[516]; 
    assign layer_0[3139] = ~(in[66] ^ in[837]); 
    assign layer_0[3140] = in[27] & ~in[808]; 
    assign layer_0[3141] = in[1000] & in[102]; 
    assign layer_0[3142] = in[431] ^ in[884]; 
    assign layer_0[3143] = ~(in[710] & in[632]); 
    assign layer_0[3144] = in[779]; 
    assign layer_0[3145] = in[918] ^ in[601]; 
    assign layer_0[3146] = in[276] & ~in[922]; 
    assign layer_0[3147] = ~(in[514] | in[608]); 
    assign layer_0[3148] = ~in[13]; 
    assign layer_0[3149] = ~in[695]; 
    assign layer_0[3150] = in[873] ^ in[837]; 
    assign layer_0[3151] = in[604]; 
    assign layer_0[3152] = ~(in[725] | in[1003]); 
    assign layer_0[3153] = ~in[160]; 
    assign layer_0[3154] = in[653] ^ in[836]; 
    assign layer_0[3155] = in[212] & ~in[482]; 
    assign layer_0[3156] = in[376] ^ in[295]; 
    assign layer_0[3157] = ~in[294]; 
    assign layer_0[3158] = ~in[836]; 
    assign layer_0[3159] = in[109] & ~in[164]; 
    assign layer_0[3160] = in[539] ^ in[603]; 
    assign layer_0[3161] = in[210]; 
    assign layer_0[3162] = ~(in[949] ^ in[952]); 
    assign layer_0[3163] = in[691] ^ in[14]; 
    assign layer_0[3164] = in[678] & in[1014]; 
    assign layer_0[3165] = ~in[881]; 
    assign layer_0[3166] = ~in[617] | (in[617] & in[664]); 
    assign layer_0[3167] = 1'b0; 
    assign layer_0[3168] = in[126] & ~in[957]; 
    assign layer_0[3169] = in[383]; 
    assign layer_0[3170] = ~in[462]; 
    assign layer_0[3171] = ~(in[47] & in[682]); 
    assign layer_0[3172] = in[41] ^ in[498]; 
    assign layer_0[3173] = ~in[249]; 
    assign layer_0[3174] = ~(in[247] ^ in[757]); 
    assign layer_0[3175] = in[931] & in[385]; 
    assign layer_0[3176] = ~in[440] | (in[648] & in[440]); 
    assign layer_0[3177] = in[919] & in[204]; 
    assign layer_0[3178] = ~in[676] | (in[955] & in[676]); 
    assign layer_0[3179] = ~(in[388] ^ in[160]); 
    assign layer_0[3180] = ~in[80] | (in[80] & in[742]); 
    assign layer_0[3181] = ~in[326]; 
    assign layer_0[3182] = in[790] ^ in[396]; 
    assign layer_0[3183] = in[36] | in[593]; 
    assign layer_0[3184] = in[555] ^ in[585]; 
    assign layer_0[3185] = in[901] ^ in[822]; 
    assign layer_0[3186] = ~(in[549] ^ in[754]); 
    assign layer_0[3187] = ~in[886] | (in[886] & in[770]); 
    assign layer_0[3188] = ~in[836] | (in[836] & in[618]); 
    assign layer_0[3189] = in[167] ^ in[372]; 
    assign layer_0[3190] = in[1014] ^ in[822]; 
    assign layer_0[3191] = ~in[147] | (in[113] & in[147]); 
    assign layer_0[3192] = in[460] ^ in[290]; 
    assign layer_0[3193] = ~(in[573] | in[996]); 
    assign layer_0[3194] = ~(in[680] & in[579]); 
    assign layer_0[3195] = ~in[902]; 
    assign layer_0[3196] = in[840] ^ in[995]; 
    assign layer_0[3197] = in[142] ^ in[467]; 
    assign layer_0[3198] = ~(in[112] ^ in[932]); 
    assign layer_0[3199] = ~in[390]; 
    assign layer_0[3200] = ~in[694]; 
    assign layer_0[3201] = in[708] ^ in[508]; 
    assign layer_0[3202] = 1'b0; 
    assign layer_0[3203] = in[9]; 
    assign layer_0[3204] = ~in[632] | (in[632] & in[775]); 
    assign layer_0[3205] = ~in[203] | (in[203] & in[638]); 
    assign layer_0[3206] = ~in[662]; 
    assign layer_0[3207] = in[344]; 
    assign layer_0[3208] = in[348] & ~in[157]; 
    assign layer_0[3209] = in[208] ^ in[454]; 
    assign layer_0[3210] = ~(in[609] | in[114]); 
    assign layer_0[3211] = in[874] ^ in[921]; 
    assign layer_0[3212] = in[556] ^ in[207]; 
    assign layer_0[3213] = ~(in[934] ^ in[933]); 
    assign layer_0[3214] = ~(in[452] ^ in[806]); 
    assign layer_0[3215] = ~in[610]; 
    assign layer_0[3216] = in[498] ^ in[751]; 
    assign layer_0[3217] = ~(in[1004] | in[419]); 
    assign layer_0[3218] = in[57]; 
    assign layer_0[3219] = in[1000] & ~in[622]; 
    assign layer_0[3220] = in[613]; 
    assign layer_0[3221] = in[520] | in[959]; 
    assign layer_0[3222] = ~in[37]; 
    assign layer_0[3223] = in[153] ^ in[42]; 
    assign layer_0[3224] = ~in[36] | (in[499] & in[36]); 
    assign layer_0[3225] = ~(in[969] & in[547]); 
    assign layer_0[3226] = in[186] & ~in[348]; 
    assign layer_0[3227] = in[564] ^ in[337]; 
    assign layer_0[3228] = in[586] & ~in[47]; 
    assign layer_0[3229] = in[490]; 
    assign layer_0[3230] = in[688] ^ in[708]; 
    assign layer_0[3231] = in[553] ^ in[599]; 
    assign layer_0[3232] = ~(in[1008] | in[942]); 
    assign layer_0[3233] = ~(in[715] ^ in[777]); 
    assign layer_0[3234] = in[235]; 
    assign layer_0[3235] = in[688] ^ in[877]; 
    assign layer_0[3236] = in[66] & in[38]; 
    assign layer_0[3237] = in[649] & ~in[286]; 
    assign layer_0[3238] = in[860] ^ in[275]; 
    assign layer_0[3239] = in[669] & ~in[849]; 
    assign layer_0[3240] = ~(in[250] & in[695]); 
    assign layer_0[3241] = in[951] ^ in[953]; 
    assign layer_0[3242] = in[125] ^ in[875]; 
    assign layer_0[3243] = in[19] ^ in[791]; 
    assign layer_0[3244] = in[418] & ~in[431]; 
    assign layer_0[3245] = in[301]; 
    assign layer_0[3246] = in[854] ^ in[905]; 
    assign layer_0[3247] = in[503] & in[983]; 
    assign layer_0[3248] = in[472] | in[440]; 
    assign layer_0[3249] = in[964]; 
    assign layer_0[3250] = ~in[147] | (in[442] & in[147]); 
    assign layer_0[3251] = ~(in[538] ^ in[532]); 
    assign layer_0[3252] = in[884] & ~in[189]; 
    assign layer_0[3253] = in[968]; 
    assign layer_0[3254] = ~(in[810] ^ in[805]); 
    assign layer_0[3255] = in[156] ^ in[35]; 
    assign layer_0[3256] = in[740] ^ in[965]; 
    assign layer_0[3257] = ~(in[277] ^ in[835]); 
    assign layer_0[3258] = in[643] & ~in[237]; 
    assign layer_0[3259] = in[491] | in[397]; 
    assign layer_0[3260] = ~(in[7] | in[925]); 
    assign layer_0[3261] = in[521] ^ in[586]; 
    assign layer_0[3262] = in[260]; 
    assign layer_0[3263] = ~in[75] | (in[75] & in[3]); 
    assign layer_0[3264] = in[750] & ~in[15]; 
    assign layer_0[3265] = ~(in[331] ^ in[252]); 
    assign layer_0[3266] = in[643] & ~in[826]; 
    assign layer_0[3267] = in[460] & ~in[68]; 
    assign layer_0[3268] = ~in[221] | (in[45] & in[221]); 
    assign layer_0[3269] = ~(in[907] ^ in[666]); 
    assign layer_0[3270] = in[37] | in[555]; 
    assign layer_0[3271] = in[250] & ~in[954]; 
    assign layer_0[3272] = ~in[555] | (in[1008] & in[555]); 
    assign layer_0[3273] = in[118] ^ in[563]; 
    assign layer_0[3274] = in[686] ^ in[933]; 
    assign layer_0[3275] = ~(in[793] | in[595]); 
    assign layer_0[3276] = ~in[476] | (in[807] & in[476]); 
    assign layer_0[3277] = ~(in[809] ^ in[667]); 
    assign layer_0[3278] = ~(in[458] | in[827]); 
    assign layer_0[3279] = ~in[460] | (in[460] & in[579]); 
    assign layer_0[3280] = in[879] ^ in[111]; 
    assign layer_0[3281] = in[699] | in[651]; 
    assign layer_0[3282] = in[657] & in[79]; 
    assign layer_0[3283] = in[840]; 
    assign layer_0[3284] = ~in[88] | (in[88] & in[81]); 
    assign layer_0[3285] = ~(in[28] & in[56]); 
    assign layer_0[3286] = ~in[964]; 
    assign layer_0[3287] = ~in[487]; 
    assign layer_0[3288] = 1'b1; 
    assign layer_0[3289] = ~(in[63] ^ in[13]); 
    assign layer_0[3290] = ~in[373]; 
    assign layer_0[3291] = ~(in[888] ^ in[65]); 
    assign layer_0[3292] = in[707] ^ in[98]; 
    assign layer_0[3293] = in[919] & ~in[603]; 
    assign layer_0[3294] = in[227] & in[615]; 
    assign layer_0[3295] = ~in[629] | (in[629] & in[700]); 
    assign layer_0[3296] = ~(in[965] | in[518]); 
    assign layer_0[3297] = ~in[476]; 
    assign layer_0[3298] = 1'b0; 
    assign layer_0[3299] = ~(in[983] ^ in[699]); 
    assign layer_0[3300] = in[920]; 
    assign layer_0[3301] = in[130] & in[686]; 
    assign layer_0[3302] = in[723]; 
    assign layer_0[3303] = in[668] ^ in[347]; 
    assign layer_0[3304] = in[715] ^ in[661]; 
    assign layer_0[3305] = in[393] & ~in[52]; 
    assign layer_0[3306] = ~in[56]; 
    assign layer_0[3307] = in[268] | in[633]; 
    assign layer_0[3308] = in[341] & ~in[671]; 
    assign layer_0[3309] = in[915] ^ in[331]; 
    assign layer_0[3310] = in[519] ^ in[307]; 
    assign layer_0[3311] = ~in[677]; 
    assign layer_0[3312] = in[835] ^ in[500]; 
    assign layer_0[3313] = ~(in[466] & in[482]); 
    assign layer_0[3314] = ~(in[364] ^ in[1017]); 
    assign layer_0[3315] = in[430] ^ in[52]; 
    assign layer_0[3316] = in[714] ^ in[672]; 
    assign layer_0[3317] = in[917]; 
    assign layer_0[3318] = ~(in[821] ^ in[288]); 
    assign layer_0[3319] = in[669] & in[860]; 
    assign layer_0[3320] = ~(in[232] & in[652]); 
    assign layer_0[3321] = ~in[587] | (in[587] & in[820]); 
    assign layer_0[3322] = in[323] ^ in[1016]; 
    assign layer_0[3323] = in[871] | in[854]; 
    assign layer_0[3324] = in[190] ^ in[490]; 
    assign layer_0[3325] = ~(in[914] ^ in[413]); 
    assign layer_0[3326] = in[921] & ~in[955]; 
    assign layer_0[3327] = in[509] ^ in[767]; 
    assign layer_0[3328] = in[745] ^ in[734]; 
    assign layer_0[3329] = in[621]; 
    assign layer_0[3330] = in[966] & in[571]; 
    assign layer_0[3331] = ~in[872]; 
    assign layer_0[3332] = ~(in[840] ^ in[889]); 
    assign layer_0[3333] = ~in[873]; 
    assign layer_0[3334] = in[584] ^ in[508]; 
    assign layer_0[3335] = ~in[446]; 
    assign layer_0[3336] = ~(in[277] & in[871]); 
    assign layer_0[3337] = in[115] & in[531]; 
    assign layer_0[3338] = ~in[385]; 
    assign layer_0[3339] = in[157] ^ in[186]; 
    assign layer_0[3340] = in[808]; 
    assign layer_0[3341] = ~(in[292] ^ in[791]); 
    assign layer_0[3342] = ~in[243]; 
    assign layer_0[3343] = 1'b0; 
    assign layer_0[3344] = ~in[37]; 
    assign layer_0[3345] = ~in[712]; 
    assign layer_0[3346] = in[59] | in[598]; 
    assign layer_0[3347] = in[944] | in[528]; 
    assign layer_0[3348] = in[857] ^ in[538]; 
    assign layer_0[3349] = ~in[193]; 
    assign layer_0[3350] = in[940] & ~in[381]; 
    assign layer_0[3351] = ~in[61]; 
    assign layer_0[3352] = ~in[148] | (in[757] & in[148]); 
    assign layer_0[3353] = in[253] | in[524]; 
    assign layer_0[3354] = 1'b0; 
    assign layer_0[3355] = in[497]; 
    assign layer_0[3356] = ~(in[102] & in[685]); 
    assign layer_0[3357] = ~(in[824] & in[431]); 
    assign layer_0[3358] = in[724] | in[397]; 
    assign layer_0[3359] = ~(in[429] ^ in[1003]); 
    assign layer_0[3360] = in[905] | in[933]; 
    assign layer_0[3361] = ~(in[100] ^ in[929]); 
    assign layer_0[3362] = in[650] | in[774]; 
    assign layer_0[3363] = ~in[394] | (in[394] & in[348]); 
    assign layer_0[3364] = in[698] ^ in[850]; 
    assign layer_0[3365] = ~in[118] | (in[267] & in[118]); 
    assign layer_0[3366] = in[789] & ~in[492]; 
    assign layer_0[3367] = ~(in[822] ^ in[696]); 
    assign layer_0[3368] = ~(in[632] & in[454]); 
    assign layer_0[3369] = in[612]; 
    assign layer_0[3370] = in[470] & ~in[793]; 
    assign layer_0[3371] = in[652] | in[405]; 
    assign layer_0[3372] = in[988] ^ in[129]; 
    assign layer_0[3373] = in[676] & in[201]; 
    assign layer_0[3374] = in[309] | in[833]; 
    assign layer_0[3375] = ~(in[518] ^ in[534]); 
    assign layer_0[3376] = in[55] & ~in[676]; 
    assign layer_0[3377] = ~in[132]; 
    assign layer_0[3378] = in[955] & ~in[898]; 
    assign layer_0[3379] = ~in[809]; 
    assign layer_0[3380] = in[317]; 
    assign layer_0[3381] = ~in[651]; 
    assign layer_0[3382] = ~in[445] | (in[445] & in[26]); 
    assign layer_0[3383] = ~(in[369] | in[39]); 
    assign layer_0[3384] = ~(in[541] ^ in[891]); 
    assign layer_0[3385] = in[603] ^ in[902]; 
    assign layer_0[3386] = ~in[137] | (in[754] & in[137]); 
    assign layer_0[3387] = in[901] ^ in[493]; 
    assign layer_0[3388] = in[131] ^ in[723]; 
    assign layer_0[3389] = ~(in[472] ^ in[819]); 
    assign layer_0[3390] = ~in[175] | (in[339] & in[175]); 
    assign layer_0[3391] = ~(in[607] ^ in[40]); 
    assign layer_0[3392] = in[905] ^ in[928]; 
    assign layer_0[3393] = ~(in[609] | in[473]); 
    assign layer_0[3394] = ~in[967]; 
    assign layer_0[3395] = ~(in[277] & in[88]); 
    assign layer_0[3396] = ~in[549]; 
    assign layer_0[3397] = in[188]; 
    assign layer_0[3398] = ~in[903] | (in[965] & in[903]); 
    assign layer_0[3399] = in[322]; 
    assign layer_0[3400] = ~(in[266] ^ in[19]); 
    assign layer_0[3401] = in[668] | in[157]; 
    assign layer_0[3402] = in[753]; 
    assign layer_0[3403] = ~in[598]; 
    assign layer_0[3404] = ~(in[72] | in[583]); 
    assign layer_0[3405] = in[984]; 
    assign layer_0[3406] = in[633] ^ in[651]; 
    assign layer_0[3407] = ~(in[353] & in[91]); 
    assign layer_0[3408] = ~in[913] | (in[308] & in[913]); 
    assign layer_0[3409] = ~(in[18] ^ in[742]); 
    assign layer_0[3410] = ~(in[682] & in[859]); 
    assign layer_0[3411] = in[763] | in[180]; 
    assign layer_0[3412] = in[917]; 
    assign layer_0[3413] = ~(in[598] | in[897]); 
    assign layer_0[3414] = in[373]; 
    assign layer_0[3415] = in[194] & ~in[799]; 
    assign layer_0[3416] = ~in[467] | (in[793] & in[467]); 
    assign layer_0[3417] = in[317] ^ in[932]; 
    assign layer_0[3418] = ~(in[968] & in[876]); 
    assign layer_0[3419] = ~(in[500] ^ in[615]); 
    assign layer_0[3420] = in[999] ^ in[506]; 
    assign layer_0[3421] = ~(in[713] ^ in[587]); 
    assign layer_0[3422] = in[8] & in[466]; 
    assign layer_0[3423] = ~in[427] | (in[427] & in[421]); 
    assign layer_0[3424] = ~(in[887] | in[586]); 
    assign layer_0[3425] = ~in[178]; 
    assign layer_0[3426] = in[63] | in[332]; 
    assign layer_0[3427] = ~in[990] | (in[609] & in[990]); 
    assign layer_0[3428] = in[110]; 
    assign layer_0[3429] = in[322] ^ in[375]; 
    assign layer_0[3430] = in[99] ^ in[641]; 
    assign layer_0[3431] = ~in[458] | (in[556] & in[458]); 
    assign layer_0[3432] = ~in[461] | (in[461] & in[18]); 
    assign layer_0[3433] = in[945] | in[18]; 
    assign layer_0[3434] = ~in[936]; 
    assign layer_0[3435] = ~(in[953] | in[715]); 
    assign layer_0[3436] = in[323] & ~in[276]; 
    assign layer_0[3437] = ~(in[275] ^ in[141]); 
    assign layer_0[3438] = ~in[62]; 
    assign layer_0[3439] = in[233] ^ in[626]; 
    assign layer_0[3440] = ~in[999] | (in[897] & in[999]); 
    assign layer_0[3441] = ~(in[418] ^ in[429]); 
    assign layer_0[3442] = in[984] ^ in[777]; 
    assign layer_0[3443] = in[680] & in[778]; 
    assign layer_0[3444] = ~(in[695] ^ in[618]); 
    assign layer_0[3445] = in[263] & ~in[379]; 
    assign layer_0[3446] = in[376] & ~in[67]; 
    assign layer_0[3447] = in[647] & ~in[764]; 
    assign layer_0[3448] = in[298] & in[826]; 
    assign layer_0[3449] = in[367] ^ in[128]; 
    assign layer_0[3450] = ~(in[936] ^ in[426]); 
    assign layer_0[3451] = in[671] | in[160]; 
    assign layer_0[3452] = ~in[47] | (in[47] & in[939]); 
    assign layer_0[3453] = in[1018] ^ in[573]; 
    assign layer_0[3454] = in[985] | in[557]; 
    assign layer_0[3455] = ~(in[133] & in[621]); 
    assign layer_0[3456] = in[227] ^ in[432]; 
    assign layer_0[3457] = in[868] & ~in[855]; 
    assign layer_0[3458] = in[673] & in[183]; 
    assign layer_0[3459] = ~in[78] | (in[78] & in[983]); 
    assign layer_0[3460] = in[404] & in[581]; 
    assign layer_0[3461] = 1'b0; 
    assign layer_0[3462] = in[3] & ~in[16]; 
    assign layer_0[3463] = in[1017] | in[638]; 
    assign layer_0[3464] = in[825] ^ in[32]; 
    assign layer_0[3465] = in[971]; 
    assign layer_0[3466] = in[906] ^ in[854]; 
    assign layer_0[3467] = ~(in[951] ^ in[875]); 
    assign layer_0[3468] = in[427] ^ in[260]; 
    assign layer_0[3469] = ~(in[62] ^ in[614]); 
    assign layer_0[3470] = in[236] ^ in[19]; 
    assign layer_0[3471] = in[760] ^ in[700]; 
    assign layer_0[3472] = ~(in[708] ^ in[276]); 
    assign layer_0[3473] = ~(in[552] ^ in[550]); 
    assign layer_0[3474] = in[243] & ~in[493]; 
    assign layer_0[3475] = in[95] & ~in[501]; 
    assign layer_0[3476] = ~in[743] | (in[743] & in[854]); 
    assign layer_0[3477] = ~(in[342] ^ in[117]); 
    assign layer_0[3478] = in[371] & ~in[888]; 
    assign layer_0[3479] = in[192] ^ in[250]; 
    assign layer_0[3480] = ~in[83] | (in[331] & in[83]); 
    assign layer_0[3481] = in[154] & in[586]; 
    assign layer_0[3482] = ~in[158] | (in[158] & in[805]); 
    assign layer_0[3483] = in[79]; 
    assign layer_0[3484] = in[832] | in[292]; 
    assign layer_0[3485] = in[1003] | in[366]; 
    assign layer_0[3486] = ~(in[855] ^ in[840]); 
    assign layer_0[3487] = ~(in[691] | in[937]); 
    assign layer_0[3488] = ~(in[937] & in[170]); 
    assign layer_0[3489] = 1'b0; 
    assign layer_0[3490] = in[169] & ~in[536]; 
    assign layer_0[3491] = in[650] ^ in[756]; 
    assign layer_0[3492] = in[411] | in[860]; 
    assign layer_0[3493] = ~in[631]; 
    assign layer_0[3494] = ~(in[202] & in[638]); 
    assign layer_0[3495] = ~in[227]; 
    assign layer_0[3496] = in[314] & in[610]; 
    assign layer_0[3497] = ~in[298] | (in[298] & in[496]); 
    assign layer_0[3498] = ~in[640]; 
    assign layer_0[3499] = in[11]; 
    assign layer_0[3500] = in[580] ^ in[371]; 
    assign layer_0[3501] = in[87] & ~in[757]; 
    assign layer_0[3502] = in[136] ^ in[46]; 
    assign layer_0[3503] = ~in[618]; 
    assign layer_0[3504] = ~(in[930] & in[624]); 
    assign layer_0[3505] = ~(in[131] ^ in[748]); 
    assign layer_0[3506] = in[205]; 
    assign layer_0[3507] = ~in[374] | (in[374] & in[871]); 
    assign layer_0[3508] = ~in[492] | (in[492] & in[597]); 
    assign layer_0[3509] = in[283] ^ in[518]; 
    assign layer_0[3510] = in[891] & ~in[498]; 
    assign layer_0[3511] = ~in[918] | (in[173] & in[918]); 
    assign layer_0[3512] = ~(in[740] ^ in[532]); 
    assign layer_0[3513] = ~(in[95] ^ in[467]); 
    assign layer_0[3514] = in[239]; 
    assign layer_0[3515] = in[935] ^ in[683]; 
    assign layer_0[3516] = ~(in[674] ^ in[866]); 
    assign layer_0[3517] = in[536] | in[254]; 
    assign layer_0[3518] = in[874] ^ in[939]; 
    assign layer_0[3519] = in[476] & in[904]; 
    assign layer_0[3520] = ~(in[175] ^ in[239]); 
    assign layer_0[3521] = ~(in[612] ^ in[604]); 
    assign layer_0[3522] = in[381] ^ in[653]; 
    assign layer_0[3523] = in[300] ^ in[291]; 
    assign layer_0[3524] = in[711] & ~in[904]; 
    assign layer_0[3525] = in[986] ^ in[620]; 
    assign layer_0[3526] = in[712] | in[855]; 
    assign layer_0[3527] = in[596] & ~in[889]; 
    assign layer_0[3528] = in[78] ^ in[728]; 
    assign layer_0[3529] = in[612] & ~in[506]; 
    assign layer_0[3530] = ~in[970]; 
    assign layer_0[3531] = ~(in[999] | in[675]); 
    assign layer_0[3532] = in[485]; 
    assign layer_0[3533] = in[35] & ~in[30]; 
    assign layer_0[3534] = ~(in[918] ^ in[867]); 
    assign layer_0[3535] = in[836] & ~in[507]; 
    assign layer_0[3536] = ~(in[850] | in[641]); 
    assign layer_0[3537] = ~(in[12] ^ in[287]); 
    assign layer_0[3538] = in[478]; 
    assign layer_0[3539] = in[195] ^ in[387]; 
    assign layer_0[3540] = 1'b0; 
    assign layer_0[3541] = ~(in[246] ^ in[956]); 
    assign layer_0[3542] = in[115] | in[100]; 
    assign layer_0[3543] = ~in[632]; 
    assign layer_0[3544] = in[7] | in[67]; 
    assign layer_0[3545] = ~(in[893] & in[201]); 
    assign layer_0[3546] = ~(in[572] | in[284]); 
    assign layer_0[3547] = in[761] ^ in[917]; 
    assign layer_0[3548] = ~in[646] | (in[646] & in[638]); 
    assign layer_0[3549] = in[874] ^ in[880]; 
    assign layer_0[3550] = in[857] | in[916]; 
    assign layer_0[3551] = in[219] & in[125]; 
    assign layer_0[3552] = ~in[910] | (in[258] & in[910]); 
    assign layer_0[3553] = ~in[667] | (in[667] & in[96]); 
    assign layer_0[3554] = in[293] ^ in[122]; 
    assign layer_0[3555] = in[885] & in[871]; 
    assign layer_0[3556] = in[916] & ~in[879]; 
    assign layer_0[3557] = in[925] & in[1001]; 
    assign layer_0[3558] = ~in[628] | (in[628] & in[478]); 
    assign layer_0[3559] = in[422] & ~in[643]; 
    assign layer_0[3560] = in[465] ^ in[211]; 
    assign layer_0[3561] = 1'b1; 
    assign layer_0[3562] = in[894] ^ in[703]; 
    assign layer_0[3563] = in[132] & in[111]; 
    assign layer_0[3564] = ~(in[843] ^ in[50]); 
    assign layer_0[3565] = 1'b0; 
    assign layer_0[3566] = ~in[718]; 
    assign layer_0[3567] = ~(in[326] | in[242]); 
    assign layer_0[3568] = in[490] ^ in[169]; 
    assign layer_0[3569] = in[607] & ~in[678]; 
    assign layer_0[3570] = in[742] | in[650]; 
    assign layer_0[3571] = ~(in[920] ^ in[721]); 
    assign layer_0[3572] = ~in[38]; 
    assign layer_0[3573] = in[433] & ~in[314]; 
    assign layer_0[3574] = ~(in[600] ^ in[66]); 
    assign layer_0[3575] = ~(in[644] ^ in[501]); 
    assign layer_0[3576] = in[621] & ~in[256]; 
    assign layer_0[3577] = ~in[185]; 
    assign layer_0[3578] = in[692] ^ in[987]; 
    assign layer_0[3579] = in[644]; 
    assign layer_0[3580] = in[504] ^ in[194]; 
    assign layer_0[3581] = ~(in[853] | in[518]); 
    assign layer_0[3582] = in[173] & ~in[32]; 
    assign layer_0[3583] = in[214] & in[670]; 
    assign layer_0[3584] = ~in[679] | (in[679] & in[301]); 
    assign layer_0[3585] = in[51] ^ in[119]; 
    assign layer_0[3586] = in[758] ^ in[595]; 
    assign layer_0[3587] = in[133] & ~in[915]; 
    assign layer_0[3588] = in[822] & in[994]; 
    assign layer_0[3589] = in[868] & ~in[501]; 
    assign layer_0[3590] = ~in[190]; 
    assign layer_0[3591] = in[657] & ~in[960]; 
    assign layer_0[3592] = ~(in[237] ^ in[163]); 
    assign layer_0[3593] = ~in[862] | (in[862] & in[222]); 
    assign layer_0[3594] = ~(in[838] ^ in[840]); 
    assign layer_0[3595] = ~(in[1014] ^ in[827]); 
    assign layer_0[3596] = in[860] ^ in[919]; 
    assign layer_0[3597] = in[676] ^ in[857]; 
    assign layer_0[3598] = ~(in[915] ^ in[568]); 
    assign layer_0[3599] = ~in[712] | (in[712] & in[757]); 
    assign layer_0[3600] = ~(in[1016] ^ in[763]); 
    assign layer_0[3601] = ~(in[969] ^ in[75]); 
    assign layer_0[3602] = in[919] & ~in[901]; 
    assign layer_0[3603] = ~(in[380] & in[823]); 
    assign layer_0[3604] = in[267] ^ in[365]; 
    assign layer_0[3605] = in[264] | in[33]; 
    assign layer_0[3606] = ~(in[300] ^ in[573]); 
    assign layer_0[3607] = in[838]; 
    assign layer_0[3608] = in[901] & ~in[986]; 
    assign layer_0[3609] = ~(in[955] | in[247]); 
    assign layer_0[3610] = ~(in[828] ^ in[923]); 
    assign layer_0[3611] = in[129] ^ in[63]; 
    assign layer_0[3612] = in[759] & in[268]; 
    assign layer_0[3613] = ~(in[731] ^ in[999]); 
    assign layer_0[3614] = in[31]; 
    assign layer_0[3615] = in[612] & ~in[877]; 
    assign layer_0[3616] = in[500] | in[676]; 
    assign layer_0[3617] = ~(in[34] | in[741]); 
    assign layer_0[3618] = 1'b0; 
    assign layer_0[3619] = in[587] & ~in[698]; 
    assign layer_0[3620] = in[98] & ~in[518]; 
    assign layer_0[3621] = in[49] | in[210]; 
    assign layer_0[3622] = in[659] ^ in[747]; 
    assign layer_0[3623] = in[450]; 
    assign layer_0[3624] = ~in[191] | (in[578] & in[191]); 
    assign layer_0[3625] = ~(in[34] | in[522]); 
    assign layer_0[3626] = in[241] ^ in[873]; 
    assign layer_0[3627] = ~(in[608] | in[1013]); 
    assign layer_0[3628] = ~in[937] | (in[872] & in[937]); 
    assign layer_0[3629] = ~(in[612] & in[926]); 
    assign layer_0[3630] = in[437] ^ in[371]; 
    assign layer_0[3631] = in[627] | in[917]; 
    assign layer_0[3632] = in[553] | in[777]; 
    assign layer_0[3633] = in[240] ^ in[119]; 
    assign layer_0[3634] = in[771] & ~in[722]; 
    assign layer_0[3635] = in[61]; 
    assign layer_0[3636] = in[468] ^ in[857]; 
    assign layer_0[3637] = ~in[424] | (in[424] & in[586]); 
    assign layer_0[3638] = ~(in[990] | in[76]); 
    assign layer_0[3639] = ~(in[194] ^ in[987]); 
    assign layer_0[3640] = ~in[38]; 
    assign layer_0[3641] = in[859] ^ in[932]; 
    assign layer_0[3642] = in[911]; 
    assign layer_0[3643] = ~(in[153] & in[457]); 
    assign layer_0[3644] = in[246] & ~in[1016]; 
    assign layer_0[3645] = ~(in[737] | in[277]); 
    assign layer_0[3646] = in[235] ^ in[175]; 
    assign layer_0[3647] = ~in[965] | (in[965] & in[919]); 
    assign layer_0[3648] = in[889] ^ in[931]; 
    assign layer_0[3649] = ~(in[623] | in[874]); 
    assign layer_0[3650] = ~(in[660] ^ in[869]); 
    assign layer_0[3651] = ~(in[43] & in[616]); 
    assign layer_0[3652] = in[56] & ~in[111]; 
    assign layer_0[3653] = in[900] & ~in[911]; 
    assign layer_0[3654] = ~in[603]; 
    assign layer_0[3655] = in[988]; 
    assign layer_0[3656] = ~in[223] | (in[828] & in[223]); 
    assign layer_0[3657] = ~(in[965] ^ in[982]); 
    assign layer_0[3658] = ~in[790]; 
    assign layer_0[3659] = in[370] & ~in[598]; 
    assign layer_0[3660] = in[842] | in[806]; 
    assign layer_0[3661] = in[727] ^ in[866]; 
    assign layer_0[3662] = ~in[115]; 
    assign layer_0[3663] = ~in[825]; 
    assign layer_0[3664] = in[623] | in[803]; 
    assign layer_0[3665] = in[774] | in[946]; 
    assign layer_0[3666] = in[853] & ~in[819]; 
    assign layer_0[3667] = in[679]; 
    assign layer_0[3668] = in[261] & in[187]; 
    assign layer_0[3669] = ~in[625] | (in[625] & in[947]); 
    assign layer_0[3670] = in[536] | in[667]; 
    assign layer_0[3671] = in[662] ^ in[520]; 
    assign layer_0[3672] = in[427] & in[489]; 
    assign layer_0[3673] = in[433] ^ in[77]; 
    assign layer_0[3674] = ~(in[1000] ^ in[809]); 
    assign layer_0[3675] = in[885] & ~in[871]; 
    assign layer_0[3676] = in[937] ^ in[982]; 
    assign layer_0[3677] = in[209] ^ in[742]; 
    assign layer_0[3678] = ~(in[694] ^ in[339]); 
    assign layer_0[3679] = ~(in[840] & in[263]); 
    assign layer_0[3680] = ~in[673] | (in[673] & in[573]); 
    assign layer_0[3681] = in[355]; 
    assign layer_0[3682] = in[403] ^ in[699]; 
    assign layer_0[3683] = ~(in[348] ^ in[621]); 
    assign layer_0[3684] = in[956] & in[133]; 
    assign layer_0[3685] = in[243] & ~in[706]; 
    assign layer_0[3686] = ~(in[793] ^ in[63]); 
    assign layer_0[3687] = ~in[947]; 
    assign layer_0[3688] = in[27] ^ in[224]; 
    assign layer_0[3689] = ~(in[11] & in[443]); 
    assign layer_0[3690] = in[516] & in[42]; 
    assign layer_0[3691] = ~in[804] | (in[246] & in[804]); 
    assign layer_0[3692] = in[328]; 
    assign layer_0[3693] = ~(in[243] ^ in[841]); 
    assign layer_0[3694] = ~in[4]; 
    assign layer_0[3695] = in[298] ^ in[748]; 
    assign layer_0[3696] = in[842] ^ in[919]; 
    assign layer_0[3697] = ~in[652] | (in[467] & in[652]); 
    assign layer_0[3698] = ~(in[684] ^ in[313]); 
    assign layer_0[3699] = ~in[262]; 
    assign layer_0[3700] = ~(in[516] | in[660]); 
    assign layer_0[3701] = ~(in[812] | in[522]); 
    assign layer_0[3702] = ~(in[756] | in[717]); 
    assign layer_0[3703] = ~(in[740] ^ in[858]); 
    assign layer_0[3704] = in[293] ^ in[538]; 
    assign layer_0[3705] = in[709] ^ in[657]; 
    assign layer_0[3706] = ~(in[300] & in[535]); 
    assign layer_0[3707] = ~(in[996] ^ in[696]); 
    assign layer_0[3708] = in[623]; 
    assign layer_0[3709] = in[30] | in[856]; 
    assign layer_0[3710] = in[479]; 
    assign layer_0[3711] = in[970] | in[30]; 
    assign layer_0[3712] = ~(in[236] & in[746]); 
    assign layer_0[3713] = in[917]; 
    assign layer_0[3714] = ~(in[666] ^ in[794]); 
    assign layer_0[3715] = ~(in[540] | in[208]); 
    assign layer_0[3716] = in[63] | in[228]; 
    assign layer_0[3717] = in[105] & ~in[973]; 
    assign layer_0[3718] = ~(in[872] | in[516]); 
    assign layer_0[3719] = in[322] & ~in[803]; 
    assign layer_0[3720] = in[1012]; 
    assign layer_0[3721] = in[921] ^ in[777]; 
    assign layer_0[3722] = in[902] ^ in[988]; 
    assign layer_0[3723] = in[555] & in[649]; 
    assign layer_0[3724] = ~(in[678] & in[447]); 
    assign layer_0[3725] = ~(in[910] ^ in[222]); 
    assign layer_0[3726] = ~(in[720] | in[611]); 
    assign layer_0[3727] = in[948] ^ in[820]; 
    assign layer_0[3728] = in[508] ^ in[519]; 
    assign layer_0[3729] = in[213] | in[930]; 
    assign layer_0[3730] = ~(in[756] | in[635]); 
    assign layer_0[3731] = ~(in[970] ^ in[969]); 
    assign layer_0[3732] = ~in[920]; 
    assign layer_0[3733] = ~(in[492] & in[876]); 
    assign layer_0[3734] = in[710]; 
    assign layer_0[3735] = in[107]; 
    assign layer_0[3736] = ~(in[968] ^ in[616]); 
    assign layer_0[3737] = ~in[80]; 
    assign layer_0[3738] = ~(in[951] ^ in[554]); 
    assign layer_0[3739] = ~in[629]; 
    assign layer_0[3740] = in[491] & in[345]; 
    assign layer_0[3741] = ~in[310]; 
    assign layer_0[3742] = ~in[969] | (in[969] & in[112]); 
    assign layer_0[3743] = in[629] ^ in[381]; 
    assign layer_0[3744] = in[672] & ~in[33]; 
    assign layer_0[3745] = 1'b0; 
    assign layer_0[3746] = in[949] ^ in[465]; 
    assign layer_0[3747] = in[705] & in[731]; 
    assign layer_0[3748] = in[362] & ~in[504]; 
    assign layer_0[3749] = in[236]; 
    assign layer_0[3750] = ~(in[161] ^ in[645]); 
    assign layer_0[3751] = in[548] ^ in[664]; 
    assign layer_0[3752] = in[82]; 
    assign layer_0[3753] = ~(in[296] | in[877]); 
    assign layer_0[3754] = ~in[267]; 
    assign layer_0[3755] = in[493] & ~in[560]; 
    assign layer_0[3756] = 1'b0; 
    assign layer_0[3757] = ~in[91]; 
    assign layer_0[3758] = ~(in[663] ^ in[590]); 
    assign layer_0[3759] = in[112] & ~in[501]; 
    assign layer_0[3760] = in[983] | in[12]; 
    assign layer_0[3761] = in[516] & ~in[349]; 
    assign layer_0[3762] = in[482] & ~in[750]; 
    assign layer_0[3763] = in[615] | in[886]; 
    assign layer_0[3764] = ~(in[819] | in[703]); 
    assign layer_0[3765] = in[567] | in[842]; 
    assign layer_0[3766] = ~(in[502] & in[550]); 
    assign layer_0[3767] = in[349] ^ in[810]; 
    assign layer_0[3768] = ~(in[633] ^ in[499]); 
    assign layer_0[3769] = ~in[917]; 
    assign layer_0[3770] = ~(in[61] & in[282]); 
    assign layer_0[3771] = in[1002] ^ in[1015]; 
    assign layer_0[3772] = in[693] ^ in[178]; 
    assign layer_0[3773] = ~(in[279] ^ in[785]); 
    assign layer_0[3774] = ~in[923] | (in[923] & in[822]); 
    assign layer_0[3775] = ~in[683] | (in[683] & in[584]); 
    assign layer_0[3776] = ~(in[86] & in[487]); 
    assign layer_0[3777] = in[300] & ~in[907]; 
    assign layer_0[3778] = in[1001] & ~in[708]; 
    assign layer_0[3779] = ~(in[50] ^ in[467]); 
    assign layer_0[3780] = ~in[374] | (in[374] & in[1021]); 
    assign layer_0[3781] = in[618] & in[348]; 
    assign layer_0[3782] = in[235] | in[499]; 
    assign layer_0[3783] = ~in[861] | (in[861] & in[245]); 
    assign layer_0[3784] = in[924] ^ in[599]; 
    assign layer_0[3785] = in[915] ^ in[363]; 
    assign layer_0[3786] = in[322] ^ in[386]; 
    assign layer_0[3787] = in[947] & ~in[657]; 
    assign layer_0[3788] = in[484] ^ in[732]; 
    assign layer_0[3789] = in[292] ^ in[372]; 
    assign layer_0[3790] = ~in[619]; 
    assign layer_0[3791] = in[471] & ~in[800]; 
    assign layer_0[3792] = in[68] ^ in[775]; 
    assign layer_0[3793] = in[311] & ~in[274]; 
    assign layer_0[3794] = in[99] & ~in[894]; 
    assign layer_0[3795] = in[79]; 
    assign layer_0[3796] = in[340] ^ in[761]; 
    assign layer_0[3797] = ~(in[247] ^ in[179]); 
    assign layer_0[3798] = ~in[531]; 
    assign layer_0[3799] = ~(in[414] & in[113]); 
    assign layer_0[3800] = ~(in[904] ^ in[890]); 
    assign layer_0[3801] = ~in[277] | (in[563] & in[277]); 
    assign layer_0[3802] = in[904]; 
    assign layer_0[3803] = ~(in[947] | in[310]); 
    assign layer_0[3804] = in[9] & ~in[643]; 
    assign layer_0[3805] = in[444] & ~in[193]; 
    assign layer_0[3806] = in[901] ^ in[970]; 
    assign layer_0[3807] = ~(in[351] | in[805]); 
    assign layer_0[3808] = ~in[979]; 
    assign layer_0[3809] = in[345] & ~in[822]; 
    assign layer_0[3810] = in[440] & in[507]; 
    assign layer_0[3811] = ~in[46] | (in[400] & in[46]); 
    assign layer_0[3812] = in[319]; 
    assign layer_0[3813] = in[986] ^ in[837]; 
    assign layer_0[3814] = in[314]; 
    assign layer_0[3815] = in[953] ^ in[384]; 
    assign layer_0[3816] = in[931] & in[466]; 
    assign layer_0[3817] = ~(in[222] | in[592]); 
    assign layer_0[3818] = ~(in[491] ^ in[745]); 
    assign layer_0[3819] = in[337]; 
    assign layer_0[3820] = ~(in[407] ^ in[611]); 
    assign layer_0[3821] = ~in[353]; 
    assign layer_0[3822] = ~in[639]; 
    assign layer_0[3823] = in[970]; 
    assign layer_0[3824] = in[13] & ~in[519]; 
    assign layer_0[3825] = ~(in[417] ^ in[497]); 
    assign layer_0[3826] = in[721] & in[968]; 
    assign layer_0[3827] = ~(in[113] ^ in[604]); 
    assign layer_0[3828] = in[373] & in[6]; 
    assign layer_0[3829] = ~(in[157] ^ in[871]); 
    assign layer_0[3830] = in[583] & ~in[974]; 
    assign layer_0[3831] = in[266] ^ in[493]; 
    assign layer_0[3832] = in[538]; 
    assign layer_0[3833] = in[677] & ~in[949]; 
    assign layer_0[3834] = ~(in[263] | in[732]); 
    assign layer_0[3835] = ~(in[941] & in[63]); 
    assign layer_0[3836] = ~in[98] | (in[98] & in[477]); 
    assign layer_0[3837] = in[267] | in[789]; 
    assign layer_0[3838] = ~in[544] | (in[544] & in[39]); 
    assign layer_0[3839] = ~(in[896] ^ in[466]); 
    assign layer_0[3840] = ~(in[189] ^ in[299]); 
    assign layer_0[3841] = ~(in[292] ^ in[626]); 
    assign layer_0[3842] = ~(in[571] | in[947]); 
    assign layer_0[3843] = ~(in[861] ^ in[818]); 
    assign layer_0[3844] = ~(in[927] & in[969]); 
    assign layer_0[3845] = in[762] | in[717]; 
    assign layer_0[3846] = in[766]; 
    assign layer_0[3847] = in[434] & in[681]; 
    assign layer_0[3848] = in[78] ^ in[744]; 
    assign layer_0[3849] = ~in[968] | (in[462] & in[968]); 
    assign layer_0[3850] = in[680] & ~in[811]; 
    assign layer_0[3851] = in[984] ^ in[774]; 
    assign layer_0[3852] = ~in[573] | (in[532] & in[573]); 
    assign layer_0[3853] = in[847] | in[266]; 
    assign layer_0[3854] = ~(in[633] ^ in[27]); 
    assign layer_0[3855] = ~in[510]; 
    assign layer_0[3856] = in[177] ^ in[468]; 
    assign layer_0[3857] = in[378]; 
    assign layer_0[3858] = in[873] | in[870]; 
    assign layer_0[3859] = in[571] & ~in[30]; 
    assign layer_0[3860] = ~(in[478] | in[890]); 
    assign layer_0[3861] = in[53] & ~in[867]; 
    assign layer_0[3862] = ~in[1018] | (in[1018] & in[754]); 
    assign layer_0[3863] = ~(in[724] ^ in[164]); 
    assign layer_0[3864] = ~in[772] | (in[872] & in[772]); 
    assign layer_0[3865] = in[640]; 
    assign layer_0[3866] = in[535] & in[694]; 
    assign layer_0[3867] = in[316] & ~in[724]; 
    assign layer_0[3868] = ~in[56] | (in[768] & in[56]); 
    assign layer_0[3869] = ~(in[84] ^ in[400]); 
    assign layer_0[3870] = ~in[607]; 
    assign layer_0[3871] = in[283] & in[1000]; 
    assign layer_0[3872] = in[916]; 
    assign layer_0[3873] = in[974] ^ in[115]; 
    assign layer_0[3874] = ~(in[85] ^ in[42]); 
    assign layer_0[3875] = ~in[931]; 
    assign layer_0[3876] = ~(in[520] ^ in[719]); 
    assign layer_0[3877] = ~in[827] | (in[477] & in[827]); 
    assign layer_0[3878] = in[812] ^ in[280]; 
    assign layer_0[3879] = in[446] ^ in[385]; 
    assign layer_0[3880] = ~in[367]; 
    assign layer_0[3881] = ~in[1001] | (in[1001] & in[554]); 
    assign layer_0[3882] = in[610] ^ in[605]; 
    assign layer_0[3883] = ~in[110]; 
    assign layer_0[3884] = ~(in[899] ^ in[729]); 
    assign layer_0[3885] = ~in[680] | (in[858] & in[680]); 
    assign layer_0[3886] = in[9] ^ in[966]; 
    assign layer_0[3887] = in[67] ^ in[458]; 
    assign layer_0[3888] = ~in[112] | (in[212] & in[112]); 
    assign layer_0[3889] = ~in[78] | (in[322] & in[78]); 
    assign layer_0[3890] = in[642] ^ in[269]; 
    assign layer_0[3891] = in[790] ^ in[938]; 
    assign layer_0[3892] = in[293] & in[760]; 
    assign layer_0[3893] = in[114] ^ in[493]; 
    assign layer_0[3894] = in[914]; 
    assign layer_0[3895] = ~in[697] | (in[697] & in[204]); 
    assign layer_0[3896] = ~(in[872] ^ in[936]); 
    assign layer_0[3897] = ~(in[31] & in[1006]); 
    assign layer_0[3898] = ~(in[682] ^ in[300]); 
    assign layer_0[3899] = ~(in[950] ^ in[853]); 
    assign layer_0[3900] = in[956] & ~in[877]; 
    assign layer_0[3901] = 1'b0; 
    assign layer_0[3902] = ~(in[428] ^ in[451]); 
    assign layer_0[3903] = ~in[396]; 
    assign layer_0[3904] = ~in[318] | (in[318] & in[821]); 
    assign layer_0[3905] = 1'b1; 
    assign layer_0[3906] = in[930] | in[30]; 
    assign layer_0[3907] = in[261] ^ in[413]; 
    assign layer_0[3908] = in[630] & ~in[172]; 
    assign layer_0[3909] = in[885]; 
    assign layer_0[3910] = in[919] ^ in[1015]; 
    assign layer_0[3911] = in[1016] ^ in[343]; 
    assign layer_0[3912] = ~in[363] | (in[363] & in[338]); 
    assign layer_0[3913] = ~in[419] | (in[419] & in[673]); 
    assign layer_0[3914] = in[468] & ~in[5]; 
    assign layer_0[3915] = ~(in[249] ^ in[946]); 
    assign layer_0[3916] = in[780]; 
    assign layer_0[3917] = ~in[964]; 
    assign layer_0[3918] = in[125] & in[200]; 
    assign layer_0[3919] = in[620]; 
    assign layer_0[3920] = in[632]; 
    assign layer_0[3921] = ~(in[219] & in[319]); 
    assign layer_0[3922] = in[915] & ~in[106]; 
    assign layer_0[3923] = in[838] ^ in[171]; 
    assign layer_0[3924] = ~in[546]; 
    assign layer_0[3925] = in[607] & ~in[739]; 
    assign layer_0[3926] = ~(in[300] ^ in[837]); 
    assign layer_0[3927] = in[428] & ~in[738]; 
    assign layer_0[3928] = ~in[35] | (in[35] & in[789]); 
    assign layer_0[3929] = in[131] ^ in[533]; 
    assign layer_0[3930] = in[853] ^ in[854]; 
    assign layer_0[3931] = in[161] ^ in[693]; 
    assign layer_0[3932] = in[966] ^ in[355]; 
    assign layer_0[3933] = ~(in[752] | in[683]); 
    assign layer_0[3934] = in[928] ^ in[197]; 
    assign layer_0[3935] = in[267] ^ in[853]; 
    assign layer_0[3936] = in[534] & ~in[19]; 
    assign layer_0[3937] = ~(in[281] | in[762]); 
    assign layer_0[3938] = ~in[74] | (in[991] & in[74]); 
    assign layer_0[3939] = ~(in[681] ^ in[662]); 
    assign layer_0[3940] = ~in[97] | (in[97] & in[707]); 
    assign layer_0[3941] = ~(in[529] | in[1002]); 
    assign layer_0[3942] = in[614] & ~in[753]; 
    assign layer_0[3943] = in[552] & ~in[468]; 
    assign layer_0[3944] = in[355] | in[12]; 
    assign layer_0[3945] = ~in[966]; 
    assign layer_0[3946] = in[555] ^ in[61]; 
    assign layer_0[3947] = in[334] & ~in[983]; 
    assign layer_0[3948] = in[986] ^ in[795]; 
    assign layer_0[3949] = in[410] ^ in[621]; 
    assign layer_0[3950] = in[10] & in[933]; 
    assign layer_0[3951] = ~(in[46] ^ in[221]); 
    assign layer_0[3952] = in[636] ^ in[988]; 
    assign layer_0[3953] = ~in[342] | (in[650] & in[342]); 
    assign layer_0[3954] = in[692]; 
    assign layer_0[3955] = ~in[517]; 
    assign layer_0[3956] = in[682] ^ in[509]; 
    assign layer_0[3957] = in[315] & ~in[508]; 
    assign layer_0[3958] = in[10] & ~in[126]; 
    assign layer_0[3959] = ~(in[891] ^ in[556]); 
    assign layer_0[3960] = in[825]; 
    assign layer_0[3961] = in[666] & in[223]; 
    assign layer_0[3962] = ~(in[643] | in[832]); 
    assign layer_0[3963] = 1'b0; 
    assign layer_0[3964] = ~(in[663] | in[986]); 
    assign layer_0[3965] = in[345] & in[697]; 
    assign layer_0[3966] = in[4]; 
    assign layer_0[3967] = in[936] & ~in[391]; 
    assign layer_0[3968] = ~(in[745] ^ in[529]); 
    assign layer_0[3969] = ~(in[641] ^ in[131]); 
    assign layer_0[3970] = ~in[387]; 
    assign layer_0[3971] = 1'b1; 
    assign layer_0[3972] = in[554] & ~in[844]; 
    assign layer_0[3973] = 1'b1; 
    assign layer_0[3974] = ~in[405]; 
    assign layer_0[3975] = in[884] & in[728]; 
    assign layer_0[3976] = ~(in[928] ^ in[93]); 
    assign layer_0[3977] = in[516] | in[794]; 
    assign layer_0[3978] = ~(in[612] | in[65]); 
    assign layer_0[3979] = in[328] ^ in[458]; 
    assign layer_0[3980] = in[930] ^ in[952]; 
    assign layer_0[3981] = ~(in[19] ^ in[822]); 
    assign layer_0[3982] = ~(in[854] ^ in[837]); 
    assign layer_0[3983] = ~in[210]; 
    assign layer_0[3984] = in[516]; 
    assign layer_0[3985] = 1'b1; 
    assign layer_0[3986] = in[147]; 
    assign layer_0[3987] = ~(in[712] ^ in[145]); 
    assign layer_0[3988] = in[639] ^ in[61]; 
    assign layer_0[3989] = ~(in[264] ^ in[859]); 
    assign layer_0[3990] = ~(in[970] ^ in[432]); 
    assign layer_0[3991] = in[758] ^ in[369]; 
    assign layer_0[3992] = in[983] | in[653]; 
    assign layer_0[3993] = ~(in[67] | in[885]); 
    assign layer_0[3994] = ~in[245]; 
    assign layer_0[3995] = in[581] ^ in[335]; 
    assign layer_0[3996] = ~(in[1011] | in[274]); 
    assign layer_0[3997] = ~in[316] | (in[316] & in[120]); 
    assign layer_0[3998] = in[1011] & in[316]; 
    assign layer_0[3999] = in[775] ^ in[791]; 
    assign layer_0[4000] = ~in[46] | (in[46] & in[605]); 
    assign layer_0[4001] = ~(in[12] ^ in[220]); 
    assign layer_0[4002] = ~in[102] | (in[86] & in[102]); 
    assign layer_0[4003] = ~(in[822] ^ in[274]); 
    assign layer_0[4004] = in[620] & ~in[627]; 
    assign layer_0[4005] = in[5] & in[868]; 
    assign layer_0[4006] = in[636] & in[221]; 
    assign layer_0[4007] = in[861]; 
    assign layer_0[4008] = ~(in[158] ^ in[267]); 
    assign layer_0[4009] = in[521]; 
    assign layer_0[4010] = in[79]; 
    assign layer_0[4011] = ~(in[615] ^ in[611]); 
    assign layer_0[4012] = ~(in[875] ^ in[904]); 
    assign layer_0[4013] = in[685] ^ in[965]; 
    assign layer_0[4014] = in[740] ^ in[412]; 
    assign layer_0[4015] = ~in[629] | (in[499] & in[629]); 
    assign layer_0[4016] = in[77] ^ in[549]; 
    assign layer_0[4017] = in[906] & ~in[581]; 
    assign layer_0[4018] = ~in[157] | (in[157] & in[813]); 
    assign layer_0[4019] = in[400] & ~in[423]; 
    assign layer_0[4020] = in[952] & ~in[604]; 
    assign layer_0[4021] = in[481] | in[639]; 
    assign layer_0[4022] = in[162] ^ in[981]; 
    assign layer_0[4023] = ~in[430] | (in[430] & in[739]); 
    assign layer_0[4024] = in[350] ^ in[835]; 
    assign layer_0[4025] = in[934] ^ in[825]; 
    assign layer_0[4026] = ~(in[871] ^ in[885]); 
    assign layer_0[4027] = in[1013] ^ in[30]; 
    assign layer_0[4028] = in[68] & ~in[262]; 
    assign layer_0[4029] = ~(in[310] ^ in[100]); 
    assign layer_0[4030] = ~(in[253] ^ in[1017]); 
    assign layer_0[4031] = ~(in[507] ^ in[268]); 
    assign layer_0[4032] = ~in[143] | (in[497] & in[143]); 
    assign layer_0[4033] = ~in[162]; 
    assign layer_0[4034] = ~in[935] | (in[935] & in[390]); 
    assign layer_0[4035] = in[612] & in[333]; 
    assign layer_0[4036] = in[695] ^ in[499]; 
    assign layer_0[4037] = in[897] & in[871]; 
    assign layer_0[4038] = in[551] & in[552]; 
    assign layer_0[4039] = in[21] & ~in[177]; 
    assign layer_0[4040] = in[614] ^ in[740]; 
    assign layer_0[4041] = ~(in[929] | in[733]); 
    assign layer_0[4042] = ~(in[868] & in[74]); 
    assign layer_0[4043] = in[315] ^ in[429]; 
    assign layer_0[4044] = ~(in[488] ^ in[255]); 
    assign layer_0[4045] = in[296] ^ in[207]; 
    assign layer_0[4046] = in[550] ^ in[677]; 
    assign layer_0[4047] = ~(in[204] | in[220]); 
    assign layer_0[4048] = in[858] & ~in[911]; 
    assign layer_0[4049] = ~(in[33] ^ in[228]); 
    assign layer_0[4050] = in[823] ^ in[842]; 
    assign layer_0[4051] = in[722]; 
    assign layer_0[4052] = in[676] ^ in[699]; 
    assign layer_0[4053] = in[253] ^ in[796]; 
    assign layer_0[4054] = ~(in[192] ^ in[318]); 
    assign layer_0[4055] = ~in[774]; 
    assign layer_0[4056] = ~(in[639] | in[47]); 
    assign layer_0[4057] = ~(in[923] ^ in[537]); 
    assign layer_0[4058] = in[917] ^ in[763]; 
    assign layer_0[4059] = ~in[706]; 
    assign layer_0[4060] = in[534] & ~in[136]; 
    assign layer_0[4061] = ~(in[690] | in[619]); 
    assign layer_0[4062] = in[1001]; 
    assign layer_0[4063] = ~in[452]; 
    assign layer_0[4064] = ~(in[857] ^ in[886]); 
    assign layer_0[4065] = ~(in[278] & in[176]); 
    assign layer_0[4066] = ~in[150]; 
    assign layer_0[4067] = in[874] & ~in[599]; 
    assign layer_0[4068] = in[469]; 
    assign layer_0[4069] = ~in[116] | (in[968] & in[116]); 
    assign layer_0[4070] = in[920]; 
    assign layer_0[4071] = in[288] ^ in[1001]; 
    assign layer_0[4072] = in[10] ^ in[922]; 
    assign layer_0[4073] = in[734] ^ in[719]; 
    assign layer_0[4074] = ~(in[130] ^ in[537]); 
    assign layer_0[4075] = in[359] & ~in[586]; 
    assign layer_0[4076] = ~(in[904] ^ in[841]); 
    assign layer_0[4077] = ~in[450]; 
    assign layer_0[4078] = in[947] & in[70]; 
    assign layer_0[4079] = in[773] | in[859]; 
    assign layer_0[4080] = ~(in[998] ^ in[100]); 
    assign layer_0[4081] = ~in[40]; 
    assign layer_0[4082] = in[948]; 
    assign layer_0[4083] = ~(in[149] ^ in[77]); 
    assign layer_0[4084] = in[871] & ~in[906]; 
    assign layer_0[4085] = in[572] ^ in[459]; 
    assign layer_0[4086] = in[21] ^ in[332]; 
    assign layer_0[4087] = ~(in[581] ^ in[428]); 
    assign layer_0[4088] = 1'b0; 
    assign layer_0[4089] = ~in[275]; 
    assign layer_0[4090] = ~in[895]; 
    assign layer_0[4091] = in[660] & in[688]; 
    assign layer_0[4092] = in[936] & in[617]; 
    assign layer_0[4093] = in[255] & ~in[222]; 
    assign layer_0[4094] = in[434] ^ in[129]; 
    assign layer_0[4095] = ~(in[906] & in[620]); 
    assign layer_0[4096] = in[985] | in[916]; 
    assign layer_0[4097] = ~in[747] | (in[300] & in[747]); 
    assign layer_0[4098] = ~(in[638] ^ in[365]); 
    assign layer_0[4099] = ~in[87]; 
    assign layer_0[4100] = ~(in[298] ^ in[997]); 
    assign layer_0[4101] = ~in[880]; 
    assign layer_0[4102] = ~in[65]; 
    assign layer_0[4103] = ~(in[638] ^ in[619]); 
    assign layer_0[4104] = in[810] ^ in[1003]; 
    assign layer_0[4105] = in[776] & in[148]; 
    assign layer_0[4106] = in[505] & ~in[553]; 
    assign layer_0[4107] = ~in[280] | (in[527] & in[280]); 
    assign layer_0[4108] = in[397]; 
    assign layer_0[4109] = ~(in[915] ^ in[571]); 
    assign layer_0[4110] = in[50] & ~in[917]; 
    assign layer_0[4111] = ~(in[771] | in[475]); 
    assign layer_0[4112] = in[95] ^ in[523]; 
    assign layer_0[4113] = in[829] | in[628]; 
    assign layer_0[4114] = ~(in[943] | in[491]); 
    assign layer_0[4115] = in[666]; 
    assign layer_0[4116] = ~(in[266] ^ in[981]); 
    assign layer_0[4117] = ~(in[382] ^ in[884]); 
    assign layer_0[4118] = in[859] ^ in[683]; 
    assign layer_0[4119] = ~in[315] | (in[464] & in[315]); 
    assign layer_0[4120] = ~(in[261] ^ in[264]); 
    assign layer_0[4121] = ~(in[711] ^ in[540]); 
    assign layer_0[4122] = in[291] & ~in[720]; 
    assign layer_0[4123] = in[331] ^ in[997]; 
    assign layer_0[4124] = ~(in[1000] ^ in[635]); 
    assign layer_0[4125] = ~(in[612] & in[603]); 
    assign layer_0[4126] = ~in[506]; 
    assign layer_0[4127] = in[103] ^ in[577]; 
    assign layer_0[4128] = ~(in[958] | in[594]); 
    assign layer_0[4129] = ~(in[826] ^ in[821]); 
    assign layer_0[4130] = ~(in[732] ^ in[822]); 
    assign layer_0[4131] = ~(in[221] | in[29]); 
    assign layer_0[4132] = in[586] | in[953]; 
    assign layer_0[4133] = in[317] ^ in[715]; 
    assign layer_0[4134] = ~(in[126] | in[637]); 
    assign layer_0[4135] = ~in[835]; 
    assign layer_0[4136] = in[731] ^ in[253]; 
    assign layer_0[4137] = in[863] ^ in[974]; 
    assign layer_0[4138] = ~(in[717] ^ in[497]); 
    assign layer_0[4139] = in[265]; 
    assign layer_0[4140] = ~(in[719] ^ in[941]); 
    assign layer_0[4141] = in[943]; 
    assign layer_0[4142] = ~(in[964] ^ in[615]); 
    assign layer_0[4143] = ~in[712] | (in[849] & in[712]); 
    assign layer_0[4144] = in[498] ^ in[209]; 
    assign layer_0[4145] = ~(in[343] | in[495]); 
    assign layer_0[4146] = 1'b1; 
    assign layer_0[4147] = ~(in[322] | in[579]); 
    assign layer_0[4148] = ~in[586] | (in[39] & in[586]); 
    assign layer_0[4149] = in[912] | in[874]; 
    assign layer_0[4150] = ~(in[446] | in[843]); 
    assign layer_0[4151] = ~in[484] | (in[484] & in[625]); 
    assign layer_0[4152] = ~(in[795] ^ in[807]); 
    assign layer_0[4153] = ~in[796] | (in[953] & in[796]); 
    assign layer_0[4154] = ~(in[520] & in[986]); 
    assign layer_0[4155] = in[142] & ~in[717]; 
    assign layer_0[4156] = 1'b0; 
    assign layer_0[4157] = ~in[711]; 
    assign layer_0[4158] = in[401]; 
    assign layer_0[4159] = in[401] & ~in[428]; 
    assign layer_0[4160] = ~(in[489] ^ in[232]); 
    assign layer_0[4161] = ~(in[878] ^ in[958]); 
    assign layer_0[4162] = ~(in[715] ^ in[81]); 
    assign layer_0[4163] = ~(in[712] | in[81]); 
    assign layer_0[4164] = in[467] ^ in[888]; 
    assign layer_0[4165] = ~(in[177] ^ in[599]); 
    assign layer_0[4166] = in[131] & ~in[613]; 
    assign layer_0[4167] = ~(in[982] ^ in[707]); 
    assign layer_0[4168] = in[952] & in[588]; 
    assign layer_0[4169] = in[618] & ~in[534]; 
    assign layer_0[4170] = in[648] ^ in[3]; 
    assign layer_0[4171] = ~(in[985] ^ in[535]); 
    assign layer_0[4172] = ~(in[938] ^ in[951]); 
    assign layer_0[4173] = in[867] & in[637]; 
    assign layer_0[4174] = ~(in[521] & in[172]); 
    assign layer_0[4175] = 1'b1; 
    assign layer_0[4176] = ~(in[890] & in[84]); 
    assign layer_0[4177] = ~in[11]; 
    assign layer_0[4178] = in[13]; 
    assign layer_0[4179] = ~in[373] | (in[1001] & in[373]); 
    assign layer_0[4180] = in[693]; 
    assign layer_0[4181] = ~in[1015] | (in[747] & in[1015]); 
    assign layer_0[4182] = in[202] ^ in[488]; 
    assign layer_0[4183] = in[45] & ~in[931]; 
    assign layer_0[4184] = in[875]; 
    assign layer_0[4185] = ~(in[175] ^ in[268]); 
    assign layer_0[4186] = ~(in[750] ^ in[730]); 
    assign layer_0[4187] = ~(in[947] | in[755]); 
    assign layer_0[4188] = in[197] & in[399]; 
    assign layer_0[4189] = in[382] & ~in[939]; 
    assign layer_0[4190] = in[855] ^ in[521]; 
    assign layer_0[4191] = ~(in[726] & in[665]); 
    assign layer_0[4192] = ~in[613] | (in[805] & in[613]); 
    assign layer_0[4193] = in[29] | in[517]; 
    assign layer_0[4194] = in[747] ^ in[938]; 
    assign layer_0[4195] = in[699]; 
    assign layer_0[4196] = in[625] | in[489]; 
    assign layer_0[4197] = in[136] & ~in[672]; 
    assign layer_0[4198] = in[253] | in[997]; 
    assign layer_0[4199] = in[477]; 
    assign layer_0[4200] = ~in[1011] | (in[1011] & in[901]); 
    assign layer_0[4201] = ~(in[792] ^ in[193]); 
    assign layer_0[4202] = ~in[716]; 
    assign layer_0[4203] = ~(in[970] & in[723]); 
    assign layer_0[4204] = ~(in[880] ^ in[276]); 
    assign layer_0[4205] = 1'b1; 
    assign layer_0[4206] = ~in[183] | (in[183] & in[160]); 
    assign layer_0[4207] = in[542] | in[905]; 
    assign layer_0[4208] = ~(in[1018] | in[597]); 
    assign layer_0[4209] = ~in[572] | (in[64] & in[572]); 
    assign layer_0[4210] = ~in[244] | (in[45] & in[244]); 
    assign layer_0[4211] = ~(in[263] | in[34]); 
    assign layer_0[4212] = in[942] & ~in[70]; 
    assign layer_0[4213] = ~(in[843] & in[709]); 
    assign layer_0[4214] = ~(in[232] ^ in[854]); 
    assign layer_0[4215] = in[278] & ~in[781]; 
    assign layer_0[4216] = in[378] & ~in[846]; 
    assign layer_0[4217] = in[887] ^ in[933]; 
    assign layer_0[4218] = ~(in[348] | in[293]); 
    assign layer_0[4219] = in[587] ^ in[970]; 
    assign layer_0[4220] = ~(in[194] ^ in[983]); 
    assign layer_0[4221] = ~(in[1013] ^ in[301]); 
    assign layer_0[4222] = ~(in[746] ^ in[897]); 
    assign layer_0[4223] = in[602] & ~in[791]; 
    assign layer_0[4224] = in[890] & ~in[785]; 
    assign layer_0[4225] = in[22]; 
    assign layer_0[4226] = in[807] | in[653]; 
    assign layer_0[4227] = ~in[630] | (in[630] & in[967]); 
    assign layer_0[4228] = in[457] ^ in[911]; 
    assign layer_0[4229] = in[665] & ~in[275]; 
    assign layer_0[4230] = in[51] & ~in[33]; 
    assign layer_0[4231] = ~(in[954] | in[483]); 
    assign layer_0[4232] = in[362] ^ in[679]; 
    assign layer_0[4233] = in[203] ^ in[425]; 
    assign layer_0[4234] = ~in[634] | (in[634] & in[723]); 
    assign layer_0[4235] = ~(in[658] & in[1016]); 
    assign layer_0[4236] = ~(in[1012] | in[852]); 
    assign layer_0[4237] = in[573] & in[420]; 
    assign layer_0[4238] = in[958] | in[65]; 
    assign layer_0[4239] = in[589] | in[632]; 
    assign layer_0[4240] = in[734] ^ in[38]; 
    assign layer_0[4241] = ~(in[697] ^ in[995]); 
    assign layer_0[4242] = ~in[918]; 
    assign layer_0[4243] = in[863] ^ in[995]; 
    assign layer_0[4244] = ~(in[253] ^ in[651]); 
    assign layer_0[4245] = 1'b1; 
    assign layer_0[4246] = ~(in[660] & in[11]); 
    assign layer_0[4247] = in[999] | in[687]; 
    assign layer_0[4248] = ~in[65]; 
    assign layer_0[4249] = in[638]; 
    assign layer_0[4250] = ~in[633] | (in[633] & in[822]); 
    assign layer_0[4251] = ~(in[192] & in[79]); 
    assign layer_0[4252] = in[173] & ~in[824]; 
    assign layer_0[4253] = in[232] & in[240]; 
    assign layer_0[4254] = ~(in[774] | in[61]); 
    assign layer_0[4255] = in[600]; 
    assign layer_0[4256] = ~in[522] | (in[522] & in[542]); 
    assign layer_0[4257] = in[476] ^ in[900]; 
    assign layer_0[4258] = in[509] & ~in[157]; 
    assign layer_0[4259] = in[582]; 
    assign layer_0[4260] = in[390] & ~in[571]; 
    assign layer_0[4261] = in[818] ^ in[637]; 
    assign layer_0[4262] = 1'b0; 
    assign layer_0[4263] = ~in[826] | (in[826] & in[808]); 
    assign layer_0[4264] = ~(in[141] | in[553]); 
    assign layer_0[4265] = 1'b1; 
    assign layer_0[4266] = 1'b1; 
    assign layer_0[4267] = ~(in[685] & in[403]); 
    assign layer_0[4268] = ~(in[955] | in[631]); 
    assign layer_0[4269] = in[569] ^ in[590]; 
    assign layer_0[4270] = in[951] & ~in[924]; 
    assign layer_0[4271] = ~(in[340] ^ in[414]); 
    assign layer_0[4272] = ~(in[589] ^ in[311]); 
    assign layer_0[4273] = ~(in[780] | in[367]); 
    assign layer_0[4274] = ~in[724]; 
    assign layer_0[4275] = in[965] & ~in[637]; 
    assign layer_0[4276] = in[22] & ~in[570]; 
    assign layer_0[4277] = ~in[587] | (in[587] & in[68]); 
    assign layer_0[4278] = ~(in[918] | in[955]); 
    assign layer_0[4279] = in[262] ^ in[759]; 
    assign layer_0[4280] = ~(in[1013] ^ in[448]); 
    assign layer_0[4281] = ~(in[657] & in[413]); 
    assign layer_0[4282] = in[461] & in[741]; 
    assign layer_0[4283] = ~(in[244] ^ in[974]); 
    assign layer_0[4284] = ~(in[728] ^ in[252]); 
    assign layer_0[4285] = ~(in[903] ^ in[996]); 
    assign layer_0[4286] = in[933]; 
    assign layer_0[4287] = in[608] ^ in[396]; 
    assign layer_0[4288] = in[759] ^ in[741]; 
    assign layer_0[4289] = in[580] & ~in[661]; 
    assign layer_0[4290] = ~in[757]; 
    assign layer_0[4291] = in[266] & in[965]; 
    assign layer_0[4292] = ~in[93] | (in[159] & in[93]); 
    assign layer_0[4293] = ~(in[82] | in[192]); 
    assign layer_0[4294] = ~(in[629] ^ in[753]); 
    assign layer_0[4295] = 1'b0; 
    assign layer_0[4296] = in[837] ^ in[29]; 
    assign layer_0[4297] = in[570] | in[128]; 
    assign layer_0[4298] = ~in[227]; 
    assign layer_0[4299] = in[965] | in[499]; 
    assign layer_0[4300] = in[919] ^ in[536]; 
    assign layer_0[4301] = in[622]; 
    assign layer_0[4302] = in[1019] & ~in[161]; 
    assign layer_0[4303] = in[603]; 
    assign layer_0[4304] = ~in[584]; 
    assign layer_0[4305] = in[709] & ~in[999]; 
    assign layer_0[4306] = ~(in[570] & in[677]); 
    assign layer_0[4307] = in[730] & in[519]; 
    assign layer_0[4308] = in[262] | in[605]; 
    assign layer_0[4309] = in[539]; 
    assign layer_0[4310] = ~(in[86] ^ in[895]); 
    assign layer_0[4311] = in[249] ^ in[240]; 
    assign layer_0[4312] = ~in[925] | (in[925] & in[720]); 
    assign layer_0[4313] = in[856] ^ in[101]; 
    assign layer_0[4314] = in[600] ^ in[953]; 
    assign layer_0[4315] = in[98] & ~in[567]; 
    assign layer_0[4316] = in[996] ^ in[246]; 
    assign layer_0[4317] = in[498]; 
    assign layer_0[4318] = in[693] ^ in[19]; 
    assign layer_0[4319] = in[91] ^ in[403]; 
    assign layer_0[4320] = in[262] & in[477]; 
    assign layer_0[4321] = in[7] & ~in[27]; 
    assign layer_0[4322] = ~(in[795] & in[298]); 
    assign layer_0[4323] = ~in[543] | (in[543] & in[526]); 
    assign layer_0[4324] = in[931]; 
    assign layer_0[4325] = ~(in[647] & in[867]); 
    assign layer_0[4326] = in[399] & ~in[38]; 
    assign layer_0[4327] = in[619]; 
    assign layer_0[4328] = in[887] | in[542]; 
    assign layer_0[4329] = ~(in[452] ^ in[806]); 
    assign layer_0[4330] = ~(in[574] ^ in[661]); 
    assign layer_0[4331] = ~(in[807] ^ in[584]); 
    assign layer_0[4332] = ~(in[715] | in[884]); 
    assign layer_0[4333] = ~in[730] | (in[730] & in[237]); 
    assign layer_0[4334] = ~(in[887] | in[461]); 
    assign layer_0[4335] = in[792] & ~in[941]; 
    assign layer_0[4336] = ~(in[22] ^ in[718]); 
    assign layer_0[4337] = in[645]; 
    assign layer_0[4338] = in[773] ^ in[162]; 
    assign layer_0[4339] = ~in[18]; 
    assign layer_0[4340] = in[371] ^ in[983]; 
    assign layer_0[4341] = ~in[534] | (in[534] & in[886]); 
    assign layer_0[4342] = ~(in[567] ^ in[199]); 
    assign layer_0[4343] = in[677] ^ in[704]; 
    assign layer_0[4344] = in[85]; 
    assign layer_0[4345] = in[221] | in[911]; 
    assign layer_0[4346] = ~(in[621] ^ in[604]); 
    assign layer_0[4347] = ~(in[682] & in[908]); 
    assign layer_0[4348] = in[148] & ~in[734]; 
    assign layer_0[4349] = in[924]; 
    assign layer_0[4350] = in[380] | in[827]; 
    assign layer_0[4351] = ~in[725] | (in[725] & in[650]); 
    assign layer_0[4352] = in[11] ^ in[659]; 
    assign layer_0[4353] = in[498]; 
    assign layer_0[4354] = in[321] & in[418]; 
    assign layer_0[4355] = ~(in[657] ^ in[8]); 
    assign layer_0[4356] = ~in[713] | (in[903] & in[713]); 
    assign layer_0[4357] = 1'b0; 
    assign layer_0[4358] = in[644] | in[764]; 
    assign layer_0[4359] = in[630] & ~in[739]; 
    assign layer_0[4360] = ~(in[578] & in[730]); 
    assign layer_0[4361] = in[997] & in[484]; 
    assign layer_0[4362] = in[952]; 
    assign layer_0[4363] = ~(in[868] ^ in[45]); 
    assign layer_0[4364] = ~(in[552] ^ in[748]); 
    assign layer_0[4365] = in[309]; 
    assign layer_0[4366] = ~(in[361] & in[759]); 
    assign layer_0[4367] = in[161] | in[355]; 
    assign layer_0[4368] = ~(in[899] & in[141]); 
    assign layer_0[4369] = in[261] & in[650]; 
    assign layer_0[4370] = ~(in[344] & in[251]); 
    assign layer_0[4371] = in[5] ^ in[263]; 
    assign layer_0[4372] = in[493]; 
    assign layer_0[4373] = ~in[36]; 
    assign layer_0[4374] = ~in[889]; 
    assign layer_0[4375] = ~(in[583] ^ in[905]); 
    assign layer_0[4376] = in[500] ^ in[95]; 
    assign layer_0[4377] = ~(in[375] & in[883]); 
    assign layer_0[4378] = ~(in[44] | in[573]); 
    assign layer_0[4379] = ~(in[777] ^ in[67]); 
    assign layer_0[4380] = ~(in[302] | in[331]); 
    assign layer_0[4381] = ~(in[180] & in[9]); 
    assign layer_0[4382] = in[12] & ~in[323]; 
    assign layer_0[4383] = ~(in[393] ^ in[476]); 
    assign layer_0[4384] = ~in[600]; 
    assign layer_0[4385] = ~in[374] | (in[491] & in[374]); 
    assign layer_0[4386] = ~in[611]; 
    assign layer_0[4387] = ~in[123] | (in[59] & in[123]); 
    assign layer_0[4388] = ~in[719]; 
    assign layer_0[4389] = in[869] ^ in[660]; 
    assign layer_0[4390] = ~in[763]; 
    assign layer_0[4391] = ~(in[882] | in[19]); 
    assign layer_0[4392] = ~(in[25] | in[618]); 
    assign layer_0[4393] = in[250] ^ in[803]; 
    assign layer_0[4394] = ~(in[206] ^ in[19]); 
    assign layer_0[4395] = ~(in[338] & in[918]); 
    assign layer_0[4396] = in[947] ^ in[183]; 
    assign layer_0[4397] = ~(in[602] ^ in[622]); 
    assign layer_0[4398] = in[604] & ~in[595]; 
    assign layer_0[4399] = ~(in[951] & in[216]); 
    assign layer_0[4400] = in[861] & ~in[209]; 
    assign layer_0[4401] = in[660] ^ in[113]; 
    assign layer_0[4402] = in[851] ^ in[627]; 
    assign layer_0[4403] = ~(in[688] & in[619]); 
    assign layer_0[4404] = in[697] & in[212]; 
    assign layer_0[4405] = in[962] | in[87]; 
    assign layer_0[4406] = in[641] ^ in[59]; 
    assign layer_0[4407] = in[111] | in[65]; 
    assign layer_0[4408] = ~in[602] | (in[360] & in[602]); 
    assign layer_0[4409] = ~in[265]; 
    assign layer_0[4410] = in[27] & ~in[745]; 
    assign layer_0[4411] = in[420] ^ in[927]; 
    assign layer_0[4412] = ~(in[179] & in[883]); 
    assign layer_0[4413] = ~in[217] | (in[217] & in[302]); 
    assign layer_0[4414] = in[238] ^ in[741]; 
    assign layer_0[4415] = ~in[595]; 
    assign layer_0[4416] = ~(in[360] & in[841]); 
    assign layer_0[4417] = ~(in[754] | in[539]); 
    assign layer_0[4418] = ~(in[938] ^ in[176]); 
    assign layer_0[4419] = ~(in[587] ^ in[839]); 
    assign layer_0[4420] = in[508] ^ in[892]; 
    assign layer_0[4421] = ~in[8] | (in[505] & in[8]); 
    assign layer_0[4422] = in[567] & ~in[533]; 
    assign layer_0[4423] = ~(in[870] ^ in[729]); 
    assign layer_0[4424] = in[758] ^ in[445]; 
    assign layer_0[4425] = ~(in[909] & in[384]); 
    assign layer_0[4426] = in[266] ^ in[276]; 
    assign layer_0[4427] = ~(in[583] ^ in[139]); 
    assign layer_0[4428] = ~(in[789] | in[100]); 
    assign layer_0[4429] = in[564] & ~in[162]; 
    assign layer_0[4430] = ~in[265]; 
    assign layer_0[4431] = ~(in[837] ^ in[755]); 
    assign layer_0[4432] = ~(in[729] ^ in[722]); 
    assign layer_0[4433] = in[42] & ~in[325]; 
    assign layer_0[4434] = ~(in[537] | in[521]); 
    assign layer_0[4435] = in[279]; 
    assign layer_0[4436] = in[906]; 
    assign layer_0[4437] = in[330] ^ in[714]; 
    assign layer_0[4438] = 1'b0; 
    assign layer_0[4439] = in[580] & in[394]; 
    assign layer_0[4440] = in[522] | in[517]; 
    assign layer_0[4441] = ~(in[623] ^ in[911]); 
    assign layer_0[4442] = ~in[583] | (in[689] & in[583]); 
    assign layer_0[4443] = in[30] ^ in[310]; 
    assign layer_0[4444] = ~(in[754] ^ in[715]); 
    assign layer_0[4445] = ~(in[601] | in[514]); 
    assign layer_0[4446] = ~in[440]; 
    assign layer_0[4447] = in[899] ^ in[719]; 
    assign layer_0[4448] = in[664]; 
    assign layer_0[4449] = ~in[615] | (in[843] & in[615]); 
    assign layer_0[4450] = ~(in[451] ^ in[322]); 
    assign layer_0[4451] = ~in[888]; 
    assign layer_0[4452] = ~(in[841] | in[827]); 
    assign layer_0[4453] = ~in[451] | (in[78] & in[451]); 
    assign layer_0[4454] = in[898] ^ in[603]; 
    assign layer_0[4455] = in[757] | in[595]; 
    assign layer_0[4456] = ~(in[728] & in[132]); 
    assign layer_0[4457] = in[397] ^ in[310]; 
    assign layer_0[4458] = in[976] | in[813]; 
    assign layer_0[4459] = ~in[502] | (in[3] & in[502]); 
    assign layer_0[4460] = in[144] & ~in[343]; 
    assign layer_0[4461] = ~in[686] | (in[686] & in[50]); 
    assign layer_0[4462] = ~(in[833] ^ in[237]); 
    assign layer_0[4463] = in[536]; 
    assign layer_0[4464] = ~in[808]; 
    assign layer_0[4465] = ~in[291]; 
    assign layer_0[4466] = in[984]; 
    assign layer_0[4467] = ~in[462] | (in[462] & in[586]); 
    assign layer_0[4468] = in[28] & in[1004]; 
    assign layer_0[4469] = in[636] & ~in[633]; 
    assign layer_0[4470] = in[174] | in[1014]; 
    assign layer_0[4471] = ~in[792] | (in[792] & in[532]); 
    assign layer_0[4472] = ~(in[936] ^ in[646]); 
    assign layer_0[4473] = in[683] & ~in[228]; 
    assign layer_0[4474] = ~in[286] | (in[286] & in[76]); 
    assign layer_0[4475] = in[565] ^ in[182]; 
    assign layer_0[4476] = in[571] ^ in[890]; 
    assign layer_0[4477] = in[601]; 
    assign layer_0[4478] = in[585] & ~in[317]; 
    assign layer_0[4479] = ~in[703] | (in[420] & in[703]); 
    assign layer_0[4480] = in[342] & in[947]; 
    assign layer_0[4481] = in[599] ^ in[924]; 
    assign layer_0[4482] = ~in[894]; 
    assign layer_0[4483] = in[788] ^ in[552]; 
    assign layer_0[4484] = ~(in[574] | in[888]); 
    assign layer_0[4485] = in[368] ^ in[928]; 
    assign layer_0[4486] = in[771] & ~in[639]; 
    assign layer_0[4487] = ~(in[594] & in[106]); 
    assign layer_0[4488] = ~(in[654] ^ in[989]); 
    assign layer_0[4489] = ~in[550] | (in[384] & in[550]); 
    assign layer_0[4490] = in[857] & ~in[225]; 
    assign layer_0[4491] = in[842] & ~in[987]; 
    assign layer_0[4492] = ~(in[193] ^ in[678]); 
    assign layer_0[4493] = ~in[598]; 
    assign layer_0[4494] = in[267]; 
    assign layer_0[4495] = in[968] ^ in[450]; 
    assign layer_0[4496] = in[347] ^ in[449]; 
    assign layer_0[4497] = in[265]; 
    assign layer_0[4498] = in[6] & ~in[793]; 
    assign layer_0[4499] = ~in[932] | (in[579] & in[932]); 
    assign layer_0[4500] = in[346] & in[245]; 
    assign layer_0[4501] = ~(in[144] | in[447]); 
    assign layer_0[4502] = ~in[253] | (in[253] & in[62]); 
    assign layer_0[4503] = in[841] & ~in[753]; 
    assign layer_0[4504] = in[418] | in[764]; 
    assign layer_0[4505] = ~(in[461] | in[177]); 
    assign layer_0[4506] = ~(in[830] & in[373]); 
    assign layer_0[4507] = in[951] & in[708]; 
    assign layer_0[4508] = ~(in[230] ^ in[536]); 
    assign layer_0[4509] = in[349]; 
    assign layer_0[4510] = ~in[699] | (in[699] & in[69]); 
    assign layer_0[4511] = in[318] | in[760]; 
    assign layer_0[4512] = ~in[825]; 
    assign layer_0[4513] = ~(in[34] ^ in[660]); 
    assign layer_0[4514] = in[360] & in[904]; 
    assign layer_0[4515] = in[998]; 
    assign layer_0[4516] = in[276] & in[699]; 
    assign layer_0[4517] = ~in[306] | (in[306] & in[827]); 
    assign layer_0[4518] = ~(in[86] | in[832]); 
    assign layer_0[4519] = ~in[765] | (in[765] & in[449]); 
    assign layer_0[4520] = in[345]; 
    assign layer_0[4521] = ~(in[571] ^ in[268]); 
    assign layer_0[4522] = ~(in[820] | in[905]); 
    assign layer_0[4523] = in[18] | in[761]; 
    assign layer_0[4524] = in[938] ^ in[59]; 
    assign layer_0[4525] = in[937] ^ in[857]; 
    assign layer_0[4526] = in[420] ^ in[580]; 
    assign layer_0[4527] = in[403] & ~in[543]; 
    assign layer_0[4528] = in[283] | in[754]; 
    assign layer_0[4529] = ~(in[206] & in[177]); 
    assign layer_0[4530] = in[568] ^ in[187]; 
    assign layer_0[4531] = ~in[611] | (in[611] & in[897]); 
    assign layer_0[4532] = ~in[490] | (in[490] & in[606]); 
    assign layer_0[4533] = in[996] ^ in[607]; 
    assign layer_0[4534] = ~in[635]; 
    assign layer_0[4535] = in[919] & ~in[583]; 
    assign layer_0[4536] = in[340]; 
    assign layer_0[4537] = in[581] ^ in[603]; 
    assign layer_0[4538] = ~(in[615] ^ in[822]); 
    assign layer_0[4539] = in[280] | in[859]; 
    assign layer_0[4540] = ~in[499] | (in[499] & in[783]); 
    assign layer_0[4541] = in[200] ^ in[189]; 
    assign layer_0[4542] = in[112]; 
    assign layer_0[4543] = ~in[871]; 
    assign layer_0[4544] = in[893] | in[739]; 
    assign layer_0[4545] = in[205] ^ in[709]; 
    assign layer_0[4546] = in[289] & ~in[296]; 
    assign layer_0[4547] = in[187] ^ in[534]; 
    assign layer_0[4548] = ~(in[29] ^ in[759]); 
    assign layer_0[4549] = ~(in[841] ^ in[742]); 
    assign layer_0[4550] = in[142] ^ in[899]; 
    assign layer_0[4551] = in[94] ^ in[261]; 
    assign layer_0[4552] = ~in[662] | (in[662] & in[536]); 
    assign layer_0[4553] = in[85] ^ in[113]; 
    assign layer_0[4554] = in[241] ^ in[942]; 
    assign layer_0[4555] = in[941] ^ in[714]; 
    assign layer_0[4556] = ~(in[809] ^ in[262]); 
    assign layer_0[4557] = 1'b0; 
    assign layer_0[4558] = in[498] | in[317]; 
    assign layer_0[4559] = ~(in[69] ^ in[932]); 
    assign layer_0[4560] = ~(in[474] ^ in[567]); 
    assign layer_0[4561] = ~(in[952] ^ in[34]); 
    assign layer_0[4562] = in[595] ^ in[954]; 
    assign layer_0[4563] = in[1002] | in[522]; 
    assign layer_0[4564] = ~in[662]; 
    assign layer_0[4565] = ~(in[588] ^ in[504]); 
    assign layer_0[4566] = in[921] ^ in[436]; 
    assign layer_0[4567] = in[900] | in[899]; 
    assign layer_0[4568] = in[579] | in[307]; 
    assign layer_0[4569] = in[689] ^ in[643]; 
    assign layer_0[4570] = in[56] & ~in[596]; 
    assign layer_0[4571] = in[87] & in[934]; 
    assign layer_0[4572] = ~(in[349] ^ in[460]); 
    assign layer_0[4573] = ~in[188] | (in[188] & in[98]); 
    assign layer_0[4574] = in[154]; 
    assign layer_0[4575] = ~(in[301] | in[450]); 
    assign layer_0[4576] = ~(in[361] ^ in[545]); 
    assign layer_0[4577] = in[532] ^ in[952]; 
    assign layer_0[4578] = ~(in[555] & in[836]); 
    assign layer_0[4579] = 1'b0; 
    assign layer_0[4580] = 1'b0; 
    assign layer_0[4581] = ~(in[701] | in[521]); 
    assign layer_0[4582] = in[725] & ~in[851]; 
    assign layer_0[4583] = ~(in[877] & in[129]); 
    assign layer_0[4584] = ~(in[737] | in[440]); 
    assign layer_0[4585] = in[858] ^ in[692]; 
    assign layer_0[4586] = in[380]; 
    assign layer_0[4587] = ~(in[353] ^ in[400]); 
    assign layer_0[4588] = ~(in[776] ^ in[860]); 
    assign layer_0[4589] = ~(in[379] | in[225]); 
    assign layer_0[4590] = ~(in[677] & in[48]); 
    assign layer_0[4591] = ~in[145] | (in[899] & in[145]); 
    assign layer_0[4592] = in[762] & ~in[335]; 
    assign layer_0[4593] = in[328] & ~in[890]; 
    assign layer_0[4594] = ~in[851]; 
    assign layer_0[4595] = ~(in[602] & in[483]); 
    assign layer_0[4596] = in[853] ^ in[874]; 
    assign layer_0[4597] = in[667] ^ in[236]; 
    assign layer_0[4598] = ~in[229] | (in[607] & in[229]); 
    assign layer_0[4599] = ~(in[971] ^ in[964]); 
    assign layer_0[4600] = ~(in[402] | in[580]); 
    assign layer_0[4601] = in[811] ^ in[673]; 
    assign layer_0[4602] = in[760] ^ in[260]; 
    assign layer_0[4603] = in[728] & ~in[142]; 
    assign layer_0[4604] = in[616] ^ in[870]; 
    assign layer_0[4605] = in[601] & in[894]; 
    assign layer_0[4606] = ~(in[329] ^ in[977]); 
    assign layer_0[4607] = ~in[395] | (in[395] & in[603]); 
    assign layer_0[4608] = ~(in[381] | in[856]); 
    assign layer_0[4609] = ~(in[506] | in[717]); 
    assign layer_0[4610] = in[716]; 
    assign layer_0[4611] = ~(in[634] | in[632]); 
    assign layer_0[4612] = ~in[967]; 
    assign layer_0[4613] = ~(in[477] ^ in[128]); 
    assign layer_0[4614] = ~(in[904] ^ in[55]); 
    assign layer_0[4615] = ~(in[373] & in[470]); 
    assign layer_0[4616] = ~in[291]; 
    assign layer_0[4617] = ~(in[698] ^ in[29]); 
    assign layer_0[4618] = in[538] ^ in[949]; 
    assign layer_0[4619] = ~in[179]; 
    assign layer_0[4620] = ~(in[763] | in[379]); 
    assign layer_0[4621] = in[841] | in[719]; 
    assign layer_0[4622] = in[462] & ~in[9]; 
    assign layer_0[4623] = ~(in[997] & in[597]); 
    assign layer_0[4624] = ~in[258] | (in[258] & in[850]); 
    assign layer_0[4625] = ~(in[875] ^ in[934]); 
    assign layer_0[4626] = ~in[878] | (in[878] & in[912]); 
    assign layer_0[4627] = ~in[301]; 
    assign layer_0[4628] = in[658]; 
    assign layer_0[4629] = ~(in[29] & in[404]); 
    assign layer_0[4630] = ~in[755]; 
    assign layer_0[4631] = ~(in[98] ^ in[666]); 
    assign layer_0[4632] = 1'b0; 
    assign layer_0[4633] = ~(in[353] & in[317]); 
    assign layer_0[4634] = ~(in[840] & in[310]); 
    assign layer_0[4635] = in[440] & ~in[780]; 
    assign layer_0[4636] = in[1002] | in[320]; 
    assign layer_0[4637] = in[492]; 
    assign layer_0[4638] = ~(in[641] | in[248]); 
    assign layer_0[4639] = ~in[615]; 
    assign layer_0[4640] = in[453] & in[45]; 
    assign layer_0[4641] = ~(in[385] ^ in[674]); 
    assign layer_0[4642] = ~(in[345] ^ in[899]); 
    assign layer_0[4643] = in[985] | in[671]; 
    assign layer_0[4644] = ~(in[282] ^ in[313]); 
    assign layer_0[4645] = in[45] ^ in[715]; 
    assign layer_0[4646] = in[352] & in[743]; 
    assign layer_0[4647] = in[619] & in[491]; 
    assign layer_0[4648] = ~in[118] | (in[477] & in[118]); 
    assign layer_0[4649] = in[101] ^ in[568]; 
    assign layer_0[4650] = ~(in[699] ^ in[76]); 
    assign layer_0[4651] = in[740] ^ in[766]; 
    assign layer_0[4652] = ~(in[191] ^ in[398]); 
    assign layer_0[4653] = ~(in[125] ^ in[420]); 
    assign layer_0[4654] = ~(in[921] ^ in[172]); 
    assign layer_0[4655] = 1'b1; 
    assign layer_0[4656] = in[504] ^ in[146]; 
    assign layer_0[4657] = ~(in[482] ^ in[492]); 
    assign layer_0[4658] = ~(in[614] ^ in[778]); 
    assign layer_0[4659] = in[983] ^ in[982]; 
    assign layer_0[4660] = in[225] ^ in[566]; 
    assign layer_0[4661] = ~in[898]; 
    assign layer_0[4662] = ~(in[597] ^ in[709]); 
    assign layer_0[4663] = in[983]; 
    assign layer_0[4664] = in[123] & ~in[936]; 
    assign layer_0[4665] = in[187] & ~in[269]; 
    assign layer_0[4666] = ~(in[551] | in[112]); 
    assign layer_0[4667] = in[981] & ~in[897]; 
    assign layer_0[4668] = ~(in[583] | in[584]); 
    assign layer_0[4669] = ~(in[333] ^ in[405]); 
    assign layer_0[4670] = in[743] ^ in[597]; 
    assign layer_0[4671] = in[469] & ~in[225]; 
    assign layer_0[4672] = in[874] & ~in[586]; 
    assign layer_0[4673] = in[210] & ~in[429]; 
    assign layer_0[4674] = ~in[396] | (in[396] & in[547]); 
    assign layer_0[4675] = ~in[493] | (in[493] & in[542]); 
    assign layer_0[4676] = ~in[591]; 
    assign layer_0[4677] = ~(in[87] | in[202]); 
    assign layer_0[4678] = ~(in[938] ^ in[553]); 
    assign layer_0[4679] = ~(in[693] & in[57]); 
    assign layer_0[4680] = in[457] & ~in[612]; 
    assign layer_0[4681] = ~in[28] | (in[28] & in[855]); 
    assign layer_0[4682] = in[239] & ~in[583]; 
    assign layer_0[4683] = ~in[986] | (in[986] & in[14]); 
    assign layer_0[4684] = in[897] & ~in[459]; 
    assign layer_0[4685] = in[858] | in[920]; 
    assign layer_0[4686] = in[291] | in[583]; 
    assign layer_0[4687] = in[842] ^ in[508]; 
    assign layer_0[4688] = ~(in[857] ^ in[262]); 
    assign layer_0[4689] = ~in[873]; 
    assign layer_0[4690] = in[923] | in[194]; 
    assign layer_0[4691] = in[258] | in[206]; 
    assign layer_0[4692] = in[256] & ~in[856]; 
    assign layer_0[4693] = in[661]; 
    assign layer_0[4694] = ~in[30] | (in[30] & in[526]); 
    assign layer_0[4695] = ~in[860]; 
    assign layer_0[4696] = in[503]; 
    assign layer_0[4697] = in[554] & ~in[980]; 
    assign layer_0[4698] = ~in[453] | (in[453] & in[980]); 
    assign layer_0[4699] = in[891] | in[144]; 
    assign layer_0[4700] = ~(in[249] ^ in[161]); 
    assign layer_0[4701] = in[70] ^ in[827]; 
    assign layer_0[4702] = ~(in[604] ^ in[735]); 
    assign layer_0[4703] = in[877] & in[378]; 
    assign layer_0[4704] = in[443]; 
    assign layer_0[4705] = ~(in[233] ^ in[939]); 
    assign layer_0[4706] = ~in[473] | (in[473] & in[239]); 
    assign layer_0[4707] = in[157] & ~in[301]; 
    assign layer_0[4708] = ~(in[381] ^ in[172]); 
    assign layer_0[4709] = in[895] ^ in[718]; 
    assign layer_0[4710] = in[184] & ~in[875]; 
    assign layer_0[4711] = in[873] & in[666]; 
    assign layer_0[4712] = in[157] | in[976]; 
    assign layer_0[4713] = in[867] ^ in[71]; 
    assign layer_0[4714] = ~in[852]; 
    assign layer_0[4715] = in[730] & ~in[923]; 
    assign layer_0[4716] = ~(in[602] ^ in[952]); 
    assign layer_0[4717] = ~in[596]; 
    assign layer_0[4718] = in[113] & ~in[886]; 
    assign layer_0[4719] = ~in[45]; 
    assign layer_0[4720] = in[209] & ~in[656]; 
    assign layer_0[4721] = in[476]; 
    assign layer_0[4722] = in[874] ^ in[983]; 
    assign layer_0[4723] = in[403] & in[239]; 
    assign layer_0[4724] = in[268] ^ in[225]; 
    assign layer_0[4725] = ~in[877] | (in[889] & in[877]); 
    assign layer_0[4726] = ~in[570]; 
    assign layer_0[4727] = in[68]; 
    assign layer_0[4728] = in[4] & ~in[14]; 
    assign layer_0[4729] = ~(in[460] ^ in[730]); 
    assign layer_0[4730] = in[489] ^ in[264]; 
    assign layer_0[4731] = in[854]; 
    assign layer_0[4732] = ~in[900] | (in[900] & in[652]); 
    assign layer_0[4733] = in[354] & ~in[269]; 
    assign layer_0[4734] = in[67] & in[343]; 
    assign layer_0[4735] = ~(in[145] ^ in[969]); 
    assign layer_0[4736] = ~(in[726] | in[948]); 
    assign layer_0[4737] = ~in[18]; 
    assign layer_0[4738] = ~in[942]; 
    assign layer_0[4739] = in[396] & in[596]; 
    assign layer_0[4740] = ~in[1015]; 
    assign layer_0[4741] = in[146] & ~in[521]; 
    assign layer_0[4742] = in[643] ^ in[233]; 
    assign layer_0[4743] = in[505] ^ in[709]; 
    assign layer_0[4744] = ~(in[254] ^ in[508]); 
    assign layer_0[4745] = ~in[420] | (in[420] & in[816]); 
    assign layer_0[4746] = ~(in[266] ^ in[1003]); 
    assign layer_0[4747] = ~(in[638] ^ in[557]); 
    assign layer_0[4748] = ~(in[35] & in[696]); 
    assign layer_0[4749] = ~(in[391] & in[238]); 
    assign layer_0[4750] = in[638] | in[610]; 
    assign layer_0[4751] = in[357]; 
    assign layer_0[4752] = in[655] & in[625]; 
    assign layer_0[4753] = ~(in[236] | in[948]); 
    assign layer_0[4754] = in[639]; 
    assign layer_0[4755] = ~in[610]; 
    assign layer_0[4756] = in[636] & in[566]; 
    assign layer_0[4757] = in[938] & ~in[80]; 
    assign layer_0[4758] = in[593] ^ in[80]; 
    assign layer_0[4759] = ~in[287]; 
    assign layer_0[4760] = ~(in[1005] & in[229]); 
    assign layer_0[4761] = ~(in[141] | in[885]); 
    assign layer_0[4762] = ~(in[698] ^ in[840]); 
    assign layer_0[4763] = ~(in[276] ^ in[520]); 
    assign layer_0[4764] = ~(in[721] ^ in[913]); 
    assign layer_0[4765] = ~(in[807] ^ in[806]); 
    assign layer_0[4766] = in[951] ^ in[651]; 
    assign layer_0[4767] = in[187] & ~in[455]; 
    assign layer_0[4768] = ~(in[791] & in[728]); 
    assign layer_0[4769] = ~in[300] | (in[872] & in[300]); 
    assign layer_0[4770] = in[655] & ~in[242]; 
    assign layer_0[4771] = in[223] & ~in[863]; 
    assign layer_0[4772] = in[967] ^ in[845]; 
    assign layer_0[4773] = in[110] ^ in[55]; 
    assign layer_0[4774] = in[618]; 
    assign layer_0[4775] = ~(in[981] ^ in[982]); 
    assign layer_0[4776] = ~(in[808] ^ in[18]); 
    assign layer_0[4777] = in[1002] & ~in[628]; 
    assign layer_0[4778] = ~in[416] | (in[26] & in[416]); 
    assign layer_0[4779] = ~(in[356] ^ in[937]); 
    assign layer_0[4780] = ~in[774] | (in[890] & in[774]); 
    assign layer_0[4781] = in[590] | in[283]; 
    assign layer_0[4782] = ~in[103] | (in[103] & in[4]); 
    assign layer_0[4783] = in[303]; 
    assign layer_0[4784] = ~in[914] | (in[593] & in[914]); 
    assign layer_0[4785] = ~(in[27] | in[852]); 
    assign layer_0[4786] = ~in[728]; 
    assign layer_0[4787] = in[633] ^ in[580]; 
    assign layer_0[4788] = ~(in[211] ^ in[890]); 
    assign layer_0[4789] = in[775] ^ in[950]; 
    assign layer_0[4790] = ~(in[660] ^ in[466]); 
    assign layer_0[4791] = ~(in[142] ^ in[499]); 
    assign layer_0[4792] = in[732] ^ in[556]; 
    assign layer_0[4793] = in[489] & in[887]; 
    assign layer_0[4794] = ~in[887] | (in[887] & in[947]); 
    assign layer_0[4795] = ~(in[267] | in[972]); 
    assign layer_0[4796] = in[55] & ~in[47]; 
    assign layer_0[4797] = ~(in[312] | in[296]); 
    assign layer_0[4798] = in[100] | in[970]; 
    assign layer_0[4799] = ~in[683] | (in[683] & in[848]); 
    assign layer_0[4800] = ~in[65] | (in[65] & in[178]); 
    assign layer_0[4801] = ~in[672]; 
    assign layer_0[4802] = ~in[680]; 
    assign layer_0[4803] = in[915] ^ in[476]; 
    assign layer_0[4804] = ~in[792]; 
    assign layer_0[4805] = in[129] | in[805]; 
    assign layer_0[4806] = ~(in[386] & in[860]); 
    assign layer_0[4807] = 1'b0; 
    assign layer_0[4808] = ~in[688] | (in[796] & in[688]); 
    assign layer_0[4809] = in[1017] ^ in[643]; 
    assign layer_0[4810] = in[25] | in[632]; 
    assign layer_0[4811] = ~in[999]; 
    assign layer_0[4812] = ~(in[1014] ^ in[483]); 
    assign layer_0[4813] = in[511] ^ in[424]; 
    assign layer_0[4814] = ~(in[139] & in[868]); 
    assign layer_0[4815] = in[744] ^ in[507]; 
    assign layer_0[4816] = ~(in[221] ^ in[876]); 
    assign layer_0[4817] = ~in[636]; 
    assign layer_0[4818] = in[931] & ~in[743]; 
    assign layer_0[4819] = in[613] & ~in[825]; 
    assign layer_0[4820] = ~(in[1005] ^ in[713]); 
    assign layer_0[4821] = in[709]; 
    assign layer_0[4822] = in[633] ^ in[910]; 
    assign layer_0[4823] = ~(in[50] ^ in[852]); 
    assign layer_0[4824] = in[981] ^ in[986]; 
    assign layer_0[4825] = ~(in[744] & in[68]); 
    assign layer_0[4826] = in[517] ^ in[568]; 
    assign layer_0[4827] = in[628] ^ in[952]; 
    assign layer_0[4828] = in[727] ^ in[995]; 
    assign layer_0[4829] = in[625] ^ in[887]; 
    assign layer_0[4830] = in[707] & in[160]; 
    assign layer_0[4831] = ~(in[296] & in[252]); 
    assign layer_0[4832] = ~(in[406] | in[48]); 
    assign layer_0[4833] = ~in[13] | (in[545] & in[13]); 
    assign layer_0[4834] = in[488] & ~in[521]; 
    assign layer_0[4835] = in[602] ^ in[945]; 
    assign layer_0[4836] = in[78] ^ in[52]; 
    assign layer_0[4837] = ~(in[633] ^ in[249]); 
    assign layer_0[4838] = ~(in[935] | in[107]); 
    assign layer_0[4839] = in[910] | in[193]; 
    assign layer_0[4840] = in[519] ^ in[275]; 
    assign layer_0[4841] = in[584] ^ in[813]; 
    assign layer_0[4842] = in[642] & in[71]; 
    assign layer_0[4843] = in[260] ^ in[710]; 
    assign layer_0[4844] = in[901] ^ in[899]; 
    assign layer_0[4845] = 1'b1; 
    assign layer_0[4846] = in[943]; 
    assign layer_0[4847] = ~in[717]; 
    assign layer_0[4848] = in[75] | in[724]; 
    assign layer_0[4849] = ~in[844] | (in[875] & in[844]); 
    assign layer_0[4850] = ~(in[886] | in[811]); 
    assign layer_0[4851] = in[838] ^ in[965]; 
    assign layer_0[4852] = in[700] & in[852]; 
    assign layer_0[4853] = in[699] & ~in[860]; 
    assign layer_0[4854] = in[912] ^ in[499]; 
    assign layer_0[4855] = ~(in[645] ^ in[984]); 
    assign layer_0[4856] = in[355] ^ in[492]; 
    assign layer_0[4857] = in[618] ^ in[511]; 
    assign layer_0[4858] = ~(in[128] ^ in[827]); 
    assign layer_0[4859] = ~(in[369] & in[672]); 
    assign layer_0[4860] = in[307] ^ in[996]; 
    assign layer_0[4861] = in[592] & in[502]; 
    assign layer_0[4862] = in[776] ^ in[596]; 
    assign layer_0[4863] = in[808] ^ in[660]; 
    assign layer_0[4864] = in[652] ^ in[260]; 
    assign layer_0[4865] = ~in[599] | (in[599] & in[857]); 
    assign layer_0[4866] = ~(in[610] | in[724]); 
    assign layer_0[4867] = in[867] | in[581]; 
    assign layer_0[4868] = in[307] & ~in[847]; 
    assign layer_0[4869] = in[254] | in[965]; 
    assign layer_0[4870] = in[859]; 
    assign layer_0[4871] = ~in[821]; 
    assign layer_0[4872] = ~in[824] | (in[824] & in[787]); 
    assign layer_0[4873] = in[552] & ~in[600]; 
    assign layer_0[4874] = in[112] & ~in[208]; 
    assign layer_0[4875] = in[419] ^ in[996]; 
    assign layer_0[4876] = in[266]; 
    assign layer_0[4877] = in[681] ^ in[221]; 
    assign layer_0[4878] = in[518]; 
    assign layer_0[4879] = in[968] ^ in[967]; 
    assign layer_0[4880] = in[635] ^ in[712]; 
    assign layer_0[4881] = in[507] ^ in[621]; 
    assign layer_0[4882] = in[326] & ~in[523]; 
    assign layer_0[4883] = ~(in[59] ^ in[980]); 
    assign layer_0[4884] = ~(in[548] ^ in[301]); 
    assign layer_0[4885] = ~(in[469] ^ in[931]); 
    assign layer_0[4886] = ~in[677] | (in[677] & in[338]); 
    assign layer_0[4887] = in[149] & in[885]; 
    assign layer_0[4888] = in[291] ^ in[999]; 
    assign layer_0[4889] = ~in[862]; 
    assign layer_0[4890] = ~(in[629] ^ in[943]); 
    assign layer_0[4891] = ~in[452]; 
    assign layer_0[4892] = in[252] & ~in[477]; 
    assign layer_0[4893] = ~in[978]; 
    assign layer_0[4894] = ~(in[609] | in[1015]); 
    assign layer_0[4895] = ~(in[366] & in[1023]); 
    assign layer_0[4896] = ~(in[955] ^ in[916]); 
    assign layer_0[4897] = in[940] ^ in[859]; 
    assign layer_0[4898] = ~(in[339] ^ in[866]); 
    assign layer_0[4899] = in[1012] | in[598]; 
    assign layer_0[4900] = in[824] & ~in[888]; 
    assign layer_0[4901] = ~(in[757] ^ in[974]); 
    assign layer_0[4902] = in[129] & ~in[614]; 
    assign layer_0[4903] = in[950] & ~in[485]; 
    assign layer_0[4904] = in[754]; 
    assign layer_0[4905] = in[632] ^ in[680]; 
    assign layer_0[4906] = ~in[267]; 
    assign layer_0[4907] = in[1001] ^ in[62]; 
    assign layer_0[4908] = in[730] & ~in[70]; 
    assign layer_0[4909] = ~(in[201] ^ in[965]); 
    assign layer_0[4910] = ~(in[354] ^ in[920]); 
    assign layer_0[4911] = ~(in[612] ^ in[824]); 
    assign layer_0[4912] = ~in[774] | (in[774] & in[968]); 
    assign layer_0[4913] = in[51]; 
    assign layer_0[4914] = ~in[702]; 
    assign layer_0[4915] = ~in[744]; 
    assign layer_0[4916] = in[715] ^ in[588]; 
    assign layer_0[4917] = ~(in[719] & in[714]); 
    assign layer_0[4918] = in[231] ^ in[907]; 
    assign layer_0[4919] = in[909]; 
    assign layer_0[4920] = ~in[952]; 
    assign layer_0[4921] = in[604]; 
    assign layer_0[4922] = in[741]; 
    assign layer_0[4923] = in[187]; 
    assign layer_0[4924] = ~(in[509] | in[877]); 
    assign layer_0[4925] = in[885] ^ in[238]; 
    assign layer_0[4926] = ~(in[673] | in[768]); 
    assign layer_0[4927] = ~(in[242] ^ in[582]); 
    assign layer_0[4928] = in[373] & ~in[260]; 
    assign layer_0[4929] = ~(in[618] ^ in[21]); 
    assign layer_0[4930] = in[919] ^ in[841]; 
    assign layer_0[4931] = ~(in[243] ^ in[788]); 
    assign layer_0[4932] = in[426] & ~in[853]; 
    assign layer_0[4933] = in[738] ^ in[4]; 
    assign layer_0[4934] = ~in[70] | (in[33] & in[70]); 
    assign layer_0[4935] = in[178] ^ in[757]; 
    assign layer_0[4936] = ~in[708]; 
    assign layer_0[4937] = ~(in[279] | in[457]); 
    assign layer_0[4938] = in[894]; 
    assign layer_0[4939] = ~in[645] | (in[645] & in[251]); 
    assign layer_0[4940] = in[811] ^ in[794]; 
    assign layer_0[4941] = in[825] & ~in[971]; 
    assign layer_0[4942] = in[262] & ~in[542]; 
    assign layer_0[4943] = ~in[4]; 
    assign layer_0[4944] = ~(in[900] ^ in[740]); 
    assign layer_0[4945] = in[443] & in[979]; 
    assign layer_0[4946] = in[145] & in[399]; 
    assign layer_0[4947] = in[553] & in[47]; 
    assign layer_0[4948] = ~(in[846] ^ in[954]); 
    assign layer_0[4949] = in[539] | in[549]; 
    assign layer_0[4950] = ~in[945] | (in[824] & in[945]); 
    assign layer_0[4951] = ~in[205] | (in[205] & in[812]); 
    assign layer_0[4952] = ~(in[112] ^ in[453]); 
    assign layer_0[4953] = ~(in[226] ^ in[999]); 
    assign layer_0[4954] = in[585] & ~in[799]; 
    assign layer_0[4955] = ~in[414] | (in[739] & in[414]); 
    assign layer_0[4956] = ~in[652]; 
    assign layer_0[4957] = ~(in[713] ^ in[840]); 
    assign layer_0[4958] = ~(in[214] ^ in[966]); 
    assign layer_0[4959] = in[564] ^ in[726]; 
    assign layer_0[4960] = in[668] ^ in[238]; 
    assign layer_0[4961] = in[680] ^ in[788]; 
    assign layer_0[4962] = in[727] ^ in[291]; 
    assign layer_0[4963] = in[549] ^ in[965]; 
    assign layer_0[4964] = in[40] & in[762]; 
    assign layer_0[4965] = in[439] & ~in[371]; 
    assign layer_0[4966] = ~(in[49] ^ in[507]); 
    assign layer_0[4967] = ~in[824] | (in[824] & in[500]); 
    assign layer_0[4968] = ~in[879]; 
    assign layer_0[4969] = ~(in[227] | in[178]); 
    assign layer_0[4970] = ~(in[821] ^ in[820]); 
    assign layer_0[4971] = in[710] & ~in[623]; 
    assign layer_0[4972] = ~in[477]; 
    assign layer_0[4973] = in[265] | in[595]; 
    assign layer_0[4974] = in[505] ^ in[933]; 
    assign layer_0[4975] = in[968] ^ in[969]; 
    assign layer_0[4976] = ~(in[807] ^ in[659]); 
    assign layer_0[4977] = ~in[996] | (in[868] & in[996]); 
    assign layer_0[4978] = in[338] | in[80]; 
    assign layer_0[4979] = in[327] & ~in[998]; 
    assign layer_0[4980] = in[538] & ~in[824]; 
    assign layer_0[4981] = in[278] ^ in[331]; 
    assign layer_0[4982] = in[688] & in[430]; 
    assign layer_0[4983] = in[327] | in[664]; 
    assign layer_0[4984] = in[565] | in[917]; 
    assign layer_0[4985] = ~in[711]; 
    assign layer_0[4986] = ~(in[749] ^ in[343]); 
    assign layer_0[4987] = in[746] & ~in[774]; 
    assign layer_0[4988] = ~(in[921] ^ in[346]); 
    assign layer_0[4989] = in[805] | in[1016]; 
    assign layer_0[4990] = in[56] & in[842]; 
    assign layer_0[4991] = ~in[611] | (in[611] & in[881]); 
    assign layer_0[4992] = ~in[206]; 
    assign layer_0[4993] = in[716] & ~in[13]; 
    assign layer_0[4994] = ~(in[129] & in[106]); 
    assign layer_0[4995] = ~in[188]; 
    assign layer_0[4996] = in[765] ^ in[810]; 
    assign layer_0[4997] = ~(in[885] ^ in[730]); 
    assign layer_0[4998] = ~in[157]; 
    assign layer_0[4999] = ~in[908] | (in[65] & in[908]); 
    assign layer_0[5000] = in[703]; 
    assign layer_0[5001] = in[712] & in[759]; 
    assign layer_0[5002] = in[653]; 
    assign layer_0[5003] = in[45] ^ in[950]; 
    assign layer_0[5004] = in[761] & ~in[433]; 
    assign layer_0[5005] = ~(in[1018] ^ in[924]); 
    assign layer_0[5006] = ~(in[627] ^ in[605]); 
    assign layer_0[5007] = in[125] | in[21]; 
    assign layer_0[5008] = ~in[196]; 
    assign layer_0[5009] = in[604] & ~in[767]; 
    assign layer_0[5010] = ~(in[153] ^ in[310]); 
    assign layer_0[5011] = ~(in[719] ^ in[888]); 
    assign layer_0[5012] = in[125] & ~in[468]; 
    assign layer_0[5013] = in[974] | in[804]; 
    assign layer_0[5014] = ~(in[98] ^ in[13]); 
    assign layer_0[5015] = in[701]; 
    assign layer_0[5016] = in[262] & in[365]; 
    assign layer_0[5017] = ~(in[116] ^ in[367]); 
    assign layer_0[5018] = ~in[858] | (in[858] & in[82]); 
    assign layer_0[5019] = ~in[728]; 
    assign layer_0[5020] = in[555]; 
    assign layer_0[5021] = ~(in[42] & in[778]); 
    assign layer_0[5022] = in[1016] | in[858]; 
    assign layer_0[5023] = ~(in[357] & in[521]); 
    assign layer_0[5024] = in[936]; 
    assign layer_0[5025] = in[835] | in[603]; 
    assign layer_0[5026] = in[935] ^ in[936]; 
    assign layer_0[5027] = in[53] ^ in[4]; 
    assign layer_0[5028] = in[334] | in[835]; 
    assign layer_0[5029] = ~in[321]; 
    assign layer_0[5030] = in[82] | in[999]; 
    assign layer_0[5031] = in[244] & ~in[858]; 
    assign layer_0[5032] = in[34] & ~in[859]; 
    assign layer_0[5033] = ~in[473] | (in[722] & in[473]); 
    assign layer_0[5034] = ~in[500] | (in[1015] & in[500]); 
    assign layer_0[5035] = ~(in[729] | in[499]); 
    assign layer_0[5036] = in[387] ^ in[414]; 
    assign layer_0[5037] = ~in[173] | (in[829] & in[173]); 
    assign layer_0[5038] = in[839] ^ in[691]; 
    assign layer_0[5039] = ~in[415]; 
    assign layer_0[5040] = in[613] ^ in[921]; 
    assign layer_0[5041] = in[598] | in[295]; 
    assign layer_0[5042] = in[859] & in[121]; 
    assign layer_0[5043] = 1'b1; 
    assign layer_0[5044] = ~(in[521] | in[284]); 
    assign layer_0[5045] = ~in[972]; 
    assign layer_0[5046] = ~in[644] | (in[644] & in[614]); 
    assign layer_0[5047] = in[625] ^ in[927]; 
    assign layer_0[5048] = ~(in[55] & in[845]); 
    assign layer_0[5049] = ~in[634] | (in[685] & in[634]); 
    assign layer_0[5050] = ~(in[980] ^ in[907]); 
    assign layer_0[5051] = 1'b1; 
    assign layer_0[5052] = ~(in[647] & in[699]); 
    assign layer_0[5053] = in[412] & in[4]; 
    assign layer_0[5054] = in[674] | in[810]; 
    assign layer_0[5055] = ~(in[914] ^ in[554]); 
    assign layer_0[5056] = ~(in[71] ^ in[857]); 
    assign layer_0[5057] = ~in[357] | (in[612] & in[357]); 
    assign layer_0[5058] = ~(in[898] & in[708]); 
    assign layer_0[5059] = ~(in[500] | in[195]); 
    assign layer_0[5060] = in[940] ^ in[853]; 
    assign layer_0[5061] = in[509]; 
    assign layer_0[5062] = ~(in[597] | in[365]); 
    assign layer_0[5063] = ~(in[325] | in[559]); 
    assign layer_0[5064] = ~in[793]; 
    assign layer_0[5065] = in[537] & ~in[501]; 
    assign layer_0[5066] = ~(in[211] | in[526]); 
    assign layer_0[5067] = in[225] ^ in[790]; 
    assign layer_0[5068] = ~(in[777] ^ in[876]); 
    assign layer_0[5069] = in[840] | in[839]; 
    assign layer_0[5070] = ~(in[544] ^ in[107]); 
    assign layer_0[5071] = ~(in[221] | in[13]); 
    assign layer_0[5072] = in[522] | in[433]; 
    assign layer_0[5073] = ~in[619] | (in[619] & in[311]); 
    assign layer_0[5074] = in[243] & ~in[177]; 
    assign layer_0[5075] = ~(in[553] & in[730]); 
    assign layer_0[5076] = ~in[858]; 
    assign layer_0[5077] = in[1015] | in[868]; 
    assign layer_0[5078] = in[499] ^ in[758]; 
    assign layer_0[5079] = ~(in[306] ^ in[500]); 
    assign layer_0[5080] = ~(in[432] & in[120]); 
    assign layer_0[5081] = in[330]; 
    assign layer_0[5082] = in[681] ^ in[699]; 
    assign layer_0[5083] = ~(in[822] & in[559]); 
    assign layer_0[5084] = ~in[236] | (in[756] & in[236]); 
    assign layer_0[5085] = in[848] & ~in[864]; 
    assign layer_0[5086] = ~(in[722] ^ in[622]); 
    assign layer_0[5087] = in[556] & in[976]; 
    assign layer_0[5088] = in[922]; 
    assign layer_0[5089] = in[350] ^ in[604]; 
    assign layer_0[5090] = in[475] | in[811]; 
    assign layer_0[5091] = ~in[572] | (in[975] & in[572]); 
    assign layer_0[5092] = in[74] | in[312]; 
    assign layer_0[5093] = in[377]; 
    assign layer_0[5094] = in[252] ^ in[744]; 
    assign layer_0[5095] = in[325] & ~in[173]; 
    assign layer_0[5096] = ~(in[689] ^ in[659]); 
    assign layer_0[5097] = in[645] ^ in[1001]; 
    assign layer_0[5098] = ~(in[760] ^ in[613]); 
    assign layer_0[5099] = in[759] | in[837]; 
    assign layer_0[5100] = ~(in[922] ^ in[583]); 
    assign layer_0[5101] = ~in[149]; 
    assign layer_0[5102] = in[324] ^ in[645]; 
    assign layer_0[5103] = in[598] ^ in[929]; 
    assign layer_0[5104] = ~(in[366] & in[398]); 
    assign layer_0[5105] = in[550] & ~in[386]; 
    assign layer_0[5106] = in[615] & in[549]; 
    assign layer_0[5107] = ~in[491]; 
    assign layer_0[5108] = ~in[924] | (in[924] & in[554]); 
    assign layer_0[5109] = ~in[518] | (in[518] & in[788]); 
    assign layer_0[5110] = ~in[479] | (in[479] & in[878]); 
    assign layer_0[5111] = in[940] ^ in[926]; 
    assign layer_0[5112] = ~(in[866] ^ in[245]); 
    assign layer_0[5113] = ~in[45] | (in[45] & in[841]); 
    assign layer_0[5114] = in[679] & in[705]; 
    assign layer_0[5115] = in[42]; 
    assign layer_0[5116] = in[157] & ~in[321]; 
    assign layer_0[5117] = in[705] ^ in[972]; 
    assign layer_0[5118] = in[451]; 
    assign layer_0[5119] = ~(in[469] ^ in[370]); 
    assign layer_0[5120] = ~(in[267] ^ in[373]); 
    assign layer_0[5121] = in[651] ^ in[600]; 
    assign layer_0[5122] = ~in[892] | (in[870] & in[892]); 
    assign layer_0[5123] = ~(in[941] ^ in[277]); 
    assign layer_0[5124] = in[350]; 
    assign layer_0[5125] = in[743] ^ in[792]; 
    assign layer_0[5126] = ~in[114]; 
    assign layer_0[5127] = in[180] ^ in[12]; 
    assign layer_0[5128] = in[968]; 
    assign layer_0[5129] = in[790]; 
    assign layer_0[5130] = in[532] ^ in[605]; 
    assign layer_0[5131] = in[532] ^ in[789]; 
    assign layer_0[5132] = in[575]; 
    assign layer_0[5133] = ~in[946]; 
    assign layer_0[5134] = ~(in[300] ^ in[291]); 
    assign layer_0[5135] = ~(in[97] ^ in[858]); 
    assign layer_0[5136] = in[803]; 
    assign layer_0[5137] = ~in[654]; 
    assign layer_0[5138] = ~(in[643] & in[657]); 
    assign layer_0[5139] = in[299] | in[955]; 
    assign layer_0[5140] = in[962] | in[565]; 
    assign layer_0[5141] = ~(in[1] ^ in[36]); 
    assign layer_0[5142] = ~in[646] | (in[646] & in[509]); 
    assign layer_0[5143] = ~in[237] | (in[141] & in[237]); 
    assign layer_0[5144] = in[661] & ~in[602]; 
    assign layer_0[5145] = ~in[46] | (in[944] & in[46]); 
    assign layer_0[5146] = ~in[927] | (in[599] & in[927]); 
    assign layer_0[5147] = ~in[440] | (in[440] & in[643]); 
    assign layer_0[5148] = in[316] & ~in[241]; 
    assign layer_0[5149] = 1'b1; 
    assign layer_0[5150] = in[971]; 
    assign layer_0[5151] = ~in[1012] | (in[825] & in[1012]); 
    assign layer_0[5152] = in[222]; 
    assign layer_0[5153] = in[1000] ^ in[234]; 
    assign layer_0[5154] = ~(in[946] ^ in[893]); 
    assign layer_0[5155] = in[242] & ~in[740]; 
    assign layer_0[5156] = ~(in[519] | in[793]); 
    assign layer_0[5157] = ~(in[305] ^ in[673]); 
    assign layer_0[5158] = ~(in[477] | in[945]); 
    assign layer_0[5159] = in[314] | in[624]; 
    assign layer_0[5160] = in[324] ^ in[537]; 
    assign layer_0[5161] = in[468] ^ in[802]; 
    assign layer_0[5162] = ~in[522]; 
    assign layer_0[5163] = ~(in[88] ^ in[456]); 
    assign layer_0[5164] = in[788] ^ in[49]; 
    assign layer_0[5165] = ~(in[322] ^ in[45]); 
    assign layer_0[5166] = in[238] ^ in[7]; 
    assign layer_0[5167] = in[911] & ~in[864]; 
    assign layer_0[5168] = ~in[840]; 
    assign layer_0[5169] = in[1015] ^ in[500]; 
    assign layer_0[5170] = ~in[58]; 
    assign layer_0[5171] = ~(in[94] ^ in[597]); 
    assign layer_0[5172] = in[550] & in[761]; 
    assign layer_0[5173] = in[664] & ~in[900]; 
    assign layer_0[5174] = in[284] ^ in[555]; 
    assign layer_0[5175] = 1'b1; 
    assign layer_0[5176] = ~in[598] | (in[598] & in[368]); 
    assign layer_0[5177] = in[454] ^ in[613]; 
    assign layer_0[5178] = ~in[170] | (in[683] & in[170]); 
    assign layer_0[5179] = in[706] ^ in[988]; 
    assign layer_0[5180] = ~(in[850] ^ in[967]); 
    assign layer_0[5181] = ~(in[746] ^ in[1000]); 
    assign layer_0[5182] = 1'b1; 
    assign layer_0[5183] = ~(in[879] ^ in[729]); 
    assign layer_0[5184] = ~in[364]; 
    assign layer_0[5185] = ~(in[222] | in[767]); 
    assign layer_0[5186] = ~(in[306] ^ in[884]); 
    assign layer_0[5187] = in[82] & in[102]; 
    assign layer_0[5188] = ~in[241]; 
    assign layer_0[5189] = in[39]; 
    assign layer_0[5190] = in[147] ^ in[707]; 
    assign layer_0[5191] = in[311] | in[568]; 
    assign layer_0[5192] = in[278] & ~in[261]; 
    assign layer_0[5193] = in[274] | in[758]; 
    assign layer_0[5194] = in[403] & ~in[125]; 
    assign layer_0[5195] = ~(in[910] & in[641]); 
    assign layer_0[5196] = in[248] ^ in[641]; 
    assign layer_0[5197] = ~in[334]; 
    assign layer_0[5198] = in[340]; 
    assign layer_0[5199] = ~(in[923] ^ in[906]); 
    assign layer_0[5200] = ~(in[937] ^ in[919]); 
    assign layer_0[5201] = in[667] ^ in[507]; 
    assign layer_0[5202] = in[19] & ~in[750]; 
    assign layer_0[5203] = ~(in[721] | in[722]); 
    assign layer_0[5204] = ~(in[1015] | in[351]); 
    assign layer_0[5205] = in[655] ^ in[55]; 
    assign layer_0[5206] = ~in[989] | (in[964] & in[989]); 
    assign layer_0[5207] = ~(in[882] ^ in[803]); 
    assign layer_0[5208] = ~in[931]; 
    assign layer_0[5209] = ~(in[709] ^ in[809]); 
    assign layer_0[5210] = ~in[1017]; 
    assign layer_0[5211] = in[732] & ~in[207]; 
    assign layer_0[5212] = in[518]; 
    assign layer_0[5213] = ~(in[637] ^ in[396]); 
    assign layer_0[5214] = ~in[797] | (in[797] & in[786]); 
    assign layer_0[5215] = ~(in[247] | in[223]); 
    assign layer_0[5216] = in[19]; 
    assign layer_0[5217] = ~in[777] | (in[777] & in[999]); 
    assign layer_0[5218] = in[829]; 
    assign layer_0[5219] = ~in[410] | (in[355] & in[410]); 
    assign layer_0[5220] = in[827] & ~in[585]; 
    assign layer_0[5221] = in[313] ^ in[262]; 
    assign layer_0[5222] = in[971]; 
    assign layer_0[5223] = ~(in[970] ^ in[12]); 
    assign layer_0[5224] = ~in[250]; 
    assign layer_0[5225] = in[808]; 
    assign layer_0[5226] = in[595]; 
    assign layer_0[5227] = in[248]; 
    assign layer_0[5228] = in[906] & ~in[228]; 
    assign layer_0[5229] = in[146] ^ in[312]; 
    assign layer_0[5230] = in[342] ^ in[182]; 
    assign layer_0[5231] = ~(in[163] | in[936]); 
    assign layer_0[5232] = ~in[430] | (in[962] & in[430]); 
    assign layer_0[5233] = in[731] & ~in[793]; 
    assign layer_0[5234] = in[141] & ~in[127]; 
    assign layer_0[5235] = ~(in[600] ^ in[726]); 
    assign layer_0[5236] = ~(in[458] ^ in[460]); 
    assign layer_0[5237] = in[599] & ~in[944]; 
    assign layer_0[5238] = in[852] & ~in[842]; 
    assign layer_0[5239] = ~(in[293] ^ in[230]); 
    assign layer_0[5240] = in[83] | in[609]; 
    assign layer_0[5241] = ~(in[760] ^ in[157]); 
    assign layer_0[5242] = in[349] & ~in[931]; 
    assign layer_0[5243] = ~in[483]; 
    assign layer_0[5244] = ~(in[160] ^ in[967]); 
    assign layer_0[5245] = ~in[868] | (in[868] & in[561]); 
    assign layer_0[5246] = ~in[297] | (in[376] & in[297]); 
    assign layer_0[5247] = in[61]; 
    assign layer_0[5248] = ~in[586]; 
    assign layer_0[5249] = in[354] ^ in[718]; 
    assign layer_0[5250] = in[453] & in[395]; 
    assign layer_0[5251] = in[154] & ~in[591]; 
    assign layer_0[5252] = in[909] ^ in[639]; 
    assign layer_0[5253] = in[964] ^ in[252]; 
    assign layer_0[5254] = ~(in[317] ^ in[924]); 
    assign layer_0[5255] = ~in[347] | (in[347] & in[837]); 
    assign layer_0[5256] = in[430] ^ in[525]; 
    assign layer_0[5257] = in[149] ^ in[415]; 
    assign layer_0[5258] = 1'b0; 
    assign layer_0[5259] = ~(in[865] | in[213]); 
    assign layer_0[5260] = ~(in[670] | in[319]); 
    assign layer_0[5261] = ~in[648] | (in[648] & in[262]); 
    assign layer_0[5262] = in[174] & ~in[434]; 
    assign layer_0[5263] = in[694] ^ in[197]; 
    assign layer_0[5264] = ~(in[291] & in[276]); 
    assign layer_0[5265] = ~in[566]; 
    assign layer_0[5266] = ~(in[741] & in[285]); 
    assign layer_0[5267] = in[700] ^ in[964]; 
    assign layer_0[5268] = ~(in[968] ^ in[961]); 
    assign layer_0[5269] = in[669] & in[626]; 
    assign layer_0[5270] = ~in[291]; 
    assign layer_0[5271] = ~in[19]; 
    assign layer_0[5272] = in[611] & in[747]; 
    assign layer_0[5273] = in[936] & ~in[891]; 
    assign layer_0[5274] = ~in[831] | (in[292] & in[831]); 
    assign layer_0[5275] = in[623] ^ in[85]; 
    assign layer_0[5276] = in[885] ^ in[646]; 
    assign layer_0[5277] = ~in[886] | (in[801] & in[886]); 
    assign layer_0[5278] = in[409]; 
    assign layer_0[5279] = in[192] & in[627]; 
    assign layer_0[5280] = in[904] & in[656]; 
    assign layer_0[5281] = in[671] | in[628]; 
    assign layer_0[5282] = in[658] ^ in[556]; 
    assign layer_0[5283] = ~in[537] | (in[537] & in[497]); 
    assign layer_0[5284] = ~in[252]; 
    assign layer_0[5285] = ~(in[980] ^ in[29]); 
    assign layer_0[5286] = ~(in[821] ^ in[662]); 
    assign layer_0[5287] = in[126]; 
    assign layer_0[5288] = ~(in[50] | in[575]); 
    assign layer_0[5289] = ~in[1015]; 
    assign layer_0[5290] = ~(in[80] | in[579]); 
    assign layer_0[5291] = 1'b1; 
    assign layer_0[5292] = in[318]; 
    assign layer_0[5293] = ~in[30]; 
    assign layer_0[5294] = in[443] & in[857]; 
    assign layer_0[5295] = ~(in[730] ^ in[496]); 
    assign layer_0[5296] = ~in[924]; 
    assign layer_0[5297] = in[524] & ~in[594]; 
    assign layer_0[5298] = ~(in[603] ^ in[584]); 
    assign layer_0[5299] = ~in[604]; 
    assign layer_0[5300] = in[380] ^ in[331]; 
    assign layer_0[5301] = in[351] & ~in[525]; 
    assign layer_0[5302] = ~in[188] | (in[188] & in[558]); 
    assign layer_0[5303] = ~(in[875] ^ in[501]); 
    assign layer_0[5304] = in[526] | in[536]; 
    assign layer_0[5305] = in[508]; 
    assign layer_0[5306] = ~in[778]; 
    assign layer_0[5307] = in[223] & ~in[730]; 
    assign layer_0[5308] = in[807]; 
    assign layer_0[5309] = ~in[419]; 
    assign layer_0[5310] = in[316] & ~in[493]; 
    assign layer_0[5311] = in[680]; 
    assign layer_0[5312] = ~(in[177] & in[664]); 
    assign layer_0[5313] = in[1017] & in[691]; 
    assign layer_0[5314] = in[822] ^ in[603]; 
    assign layer_0[5315] = 1'b0; 
    assign layer_0[5316] = in[982] & ~in[956]; 
    assign layer_0[5317] = ~(in[906] | in[27]); 
    assign layer_0[5318] = in[466] ^ in[61]; 
    assign layer_0[5319] = ~(in[904] | in[178]); 
    assign layer_0[5320] = ~in[648]; 
    assign layer_0[5321] = in[334] & in[645]; 
    assign layer_0[5322] = ~in[59] | (in[516] & in[59]); 
    assign layer_0[5323] = ~in[654]; 
    assign layer_0[5324] = in[587] & in[340]; 
    assign layer_0[5325] = ~(in[679] ^ in[774]); 
    assign layer_0[5326] = in[177] ^ in[931]; 
    assign layer_0[5327] = ~(in[983] ^ in[163]); 
    assign layer_0[5328] = in[650] & ~in[989]; 
    assign layer_0[5329] = in[697] | in[978]; 
    assign layer_0[5330] = ~in[872]; 
    assign layer_0[5331] = in[478]; 
    assign layer_0[5332] = in[867] & in[859]; 
    assign layer_0[5333] = ~(in[301] ^ in[927]); 
    assign layer_0[5334] = in[264]; 
    assign layer_0[5335] = ~(in[650] ^ in[795]); 
    assign layer_0[5336] = ~in[630]; 
    assign layer_0[5337] = ~(in[1006] ^ in[582]); 
    assign layer_0[5338] = ~in[614] | (in[614] & in[160]); 
    assign layer_0[5339] = 1'b0; 
    assign layer_0[5340] = ~(in[143] ^ in[8]); 
    assign layer_0[5341] = in[176] | in[241]; 
    assign layer_0[5342] = ~(in[411] ^ in[84]); 
    assign layer_0[5343] = ~(in[538] ^ in[500]); 
    assign layer_0[5344] = ~in[301]; 
    assign layer_0[5345] = in[926] & ~in[67]; 
    assign layer_0[5346] = in[731] ^ in[428]; 
    assign layer_0[5347] = ~in[74] | (in[714] & in[74]); 
    assign layer_0[5348] = ~in[118] | (in[644] & in[118]); 
    assign layer_0[5349] = in[804] ^ in[184]; 
    assign layer_0[5350] = in[806]; 
    assign layer_0[5351] = ~in[955]; 
    assign layer_0[5352] = in[290] & ~in[28]; 
    assign layer_0[5353] = in[597] & in[491]; 
    assign layer_0[5354] = in[204] | in[402]; 
    assign layer_0[5355] = ~(in[871] & in[523]); 
    assign layer_0[5356] = ~(in[98] ^ in[493]); 
    assign layer_0[5357] = ~in[448]; 
    assign layer_0[5358] = ~(in[721] & in[661]); 
    assign layer_0[5359] = ~(in[949] ^ in[483]); 
    assign layer_0[5360] = ~(in[68] | in[899]); 
    assign layer_0[5361] = ~(in[821] & in[762]); 
    assign layer_0[5362] = in[550] & ~in[902]; 
    assign layer_0[5363] = ~in[791] | (in[842] & in[791]); 
    assign layer_0[5364] = ~in[91] | (in[91] & in[156]); 
    assign layer_0[5365] = ~(in[331] ^ in[618]); 
    assign layer_0[5366] = in[630] ^ in[972]; 
    assign layer_0[5367] = ~in[488] | (in[488] & in[509]); 
    assign layer_0[5368] = ~in[434]; 
    assign layer_0[5369] = ~(in[105] ^ in[300]); 
    assign layer_0[5370] = ~(in[19] ^ in[569]); 
    assign layer_0[5371] = in[263]; 
    assign layer_0[5372] = ~in[365] | (in[769] & in[365]); 
    assign layer_0[5373] = ~(in[276] ^ in[83]); 
    assign layer_0[5374] = ~(in[518] ^ in[969]); 
    assign layer_0[5375] = ~(in[925] ^ in[905]); 
    assign layer_0[5376] = in[143]; 
    assign layer_0[5377] = in[918] ^ in[934]; 
    assign layer_0[5378] = ~(in[1001] ^ in[1000]); 
    assign layer_0[5379] = in[921]; 
    assign layer_0[5380] = in[110]; 
    assign layer_0[5381] = ~(in[780] | in[545]); 
    assign layer_0[5382] = ~in[947] | (in[240] & in[947]); 
    assign layer_0[5383] = in[724]; 
    assign layer_0[5384] = 1'b0; 
    assign layer_0[5385] = in[810] & ~in[841]; 
    assign layer_0[5386] = in[345]; 
    assign layer_0[5387] = ~in[254]; 
    assign layer_0[5388] = in[717] & ~in[616]; 
    assign layer_0[5389] = in[879] ^ in[167]; 
    assign layer_0[5390] = ~in[947] | (in[947] & in[4]); 
    assign layer_0[5391] = ~in[47] | (in[47] & in[615]); 
    assign layer_0[5392] = ~in[563]; 
    assign layer_0[5393] = ~(in[309] ^ in[900]); 
    assign layer_0[5394] = in[792] ^ in[922]; 
    assign layer_0[5395] = in[808] ^ in[792]; 
    assign layer_0[5396] = in[229] ^ in[210]; 
    assign layer_0[5397] = ~(in[21] & in[253]); 
    assign layer_0[5398] = ~(in[264] & in[265]); 
    assign layer_0[5399] = in[948] & in[666]; 
    assign layer_0[5400] = in[655] & ~in[790]; 
    assign layer_0[5401] = in[712] ^ in[452]; 
    assign layer_0[5402] = in[244] ^ in[575]; 
    assign layer_0[5403] = ~in[665] | (in[665] & in[635]); 
    assign layer_0[5404] = in[914] ^ in[625]; 
    assign layer_0[5405] = in[234] & ~in[2]; 
    assign layer_0[5406] = in[221] & ~in[837]; 
    assign layer_0[5407] = ~in[795]; 
    assign layer_0[5408] = ~in[467]; 
    assign layer_0[5409] = in[822] ^ in[697]; 
    assign layer_0[5410] = ~in[894]; 
    assign layer_0[5411] = in[777] ^ in[174]; 
    assign layer_0[5412] = ~(in[382] ^ in[94]); 
    assign layer_0[5413] = ~(in[74] & in[633]); 
    assign layer_0[5414] = ~(in[759] ^ in[555]); 
    assign layer_0[5415] = ~(in[267] | in[810]); 
    assign layer_0[5416] = in[17]; 
    assign layer_0[5417] = ~(in[641] ^ in[938]); 
    assign layer_0[5418] = ~(in[861] | in[640]); 
    assign layer_0[5419] = ~(in[654] ^ in[605]); 
    assign layer_0[5420] = ~(in[530] | in[690]); 
    assign layer_0[5421] = ~in[341] | (in[341] & in[768]); 
    assign layer_0[5422] = ~in[926] | (in[926] & in[729]); 
    assign layer_0[5423] = in[381] ^ in[817]; 
    assign layer_0[5424] = in[92]; 
    assign layer_0[5425] = ~in[470] | (in[892] & in[470]); 
    assign layer_0[5426] = in[598] | in[971]; 
    assign layer_0[5427] = in[13] & in[180]; 
    assign layer_0[5428] = in[242] & ~in[52]; 
    assign layer_0[5429] = in[1012] | in[700]; 
    assign layer_0[5430] = ~(in[300] ^ in[731]); 
    assign layer_0[5431] = in[983] ^ in[314]; 
    assign layer_0[5432] = ~in[619] | (in[619] & in[591]); 
    assign layer_0[5433] = in[50] | in[447]; 
    assign layer_0[5434] = ~in[620] | (in[620] & in[995]); 
    assign layer_0[5435] = in[65] | in[729]; 
    assign layer_0[5436] = ~(in[886] | in[688]); 
    assign layer_0[5437] = ~in[632] | (in[578] & in[632]); 
    assign layer_0[5438] = ~in[629]; 
    assign layer_0[5439] = in[475] ^ in[647]; 
    assign layer_0[5440] = ~in[433] | (in[266] & in[433]); 
    assign layer_0[5441] = ~in[100] | (in[986] & in[100]); 
    assign layer_0[5442] = ~(in[366] ^ in[995]); 
    assign layer_0[5443] = in[60] & ~in[275]; 
    assign layer_0[5444] = ~in[221] | (in[221] & in[748]); 
    assign layer_0[5445] = ~in[639] | (in[639] & in[597]); 
    assign layer_0[5446] = in[714]; 
    assign layer_0[5447] = in[583] & ~in[286]; 
    assign layer_0[5448] = in[967] ^ in[612]; 
    assign layer_0[5449] = in[195] & ~in[970]; 
    assign layer_0[5450] = ~(in[351] ^ in[103]); 
    assign layer_0[5451] = in[671] & ~in[45]; 
    assign layer_0[5452] = ~(in[561] | in[68]); 
    assign layer_0[5453] = in[135] & ~in[780]; 
    assign layer_0[5454] = in[493] & in[489]; 
    assign layer_0[5455] = in[460] ^ in[275]; 
    assign layer_0[5456] = ~in[373]; 
    assign layer_0[5457] = in[261] ^ in[276]; 
    assign layer_0[5458] = ~in[599] | (in[621] & in[599]); 
    assign layer_0[5459] = ~in[500]; 
    assign layer_0[5460] = in[68] ^ in[941]; 
    assign layer_0[5461] = ~(in[49] ^ in[872]); 
    assign layer_0[5462] = ~(in[872] ^ in[568]); 
    assign layer_0[5463] = in[915] ^ in[912]; 
    assign layer_0[5464] = in[280]; 
    assign layer_0[5465] = ~in[539]; 
    assign layer_0[5466] = in[596] & ~in[462]; 
    assign layer_0[5467] = ~(in[310] | in[704]); 
    assign layer_0[5468] = ~(in[695] | in[664]); 
    assign layer_0[5469] = in[214] | in[37]; 
    assign layer_0[5470] = in[967] & ~in[763]; 
    assign layer_0[5471] = 1'b0; 
    assign layer_0[5472] = ~(in[147] ^ in[456]); 
    assign layer_0[5473] = in[94] | in[891]; 
    assign layer_0[5474] = 1'b1; 
    assign layer_0[5475] = ~in[428] | (in[428] & in[734]); 
    assign layer_0[5476] = 1'b1; 
    assign layer_0[5477] = ~in[948]; 
    assign layer_0[5478] = 1'b0; 
    assign layer_0[5479] = ~(in[209] ^ in[29]); 
    assign layer_0[5480] = ~in[767] | (in[368] & in[767]); 
    assign layer_0[5481] = in[487] | in[917]; 
    assign layer_0[5482] = ~in[760] | (in[760] & in[600]); 
    assign layer_0[5483] = in[774] | in[951]; 
    assign layer_0[5484] = in[631] ^ in[757]; 
    assign layer_0[5485] = in[461] ^ in[481]; 
    assign layer_0[5486] = in[46] ^ in[207]; 
    assign layer_0[5487] = in[62] | in[1013]; 
    assign layer_0[5488] = ~in[614] | (in[656] & in[614]); 
    assign layer_0[5489] = ~in[65] | (in[65] & in[401]); 
    assign layer_0[5490] = ~in[448] | (in[221] & in[448]); 
    assign layer_0[5491] = in[659] & in[665]; 
    assign layer_0[5492] = in[984] ^ in[835]; 
    assign layer_0[5493] = in[484] ^ in[386]; 
    assign layer_0[5494] = ~(in[679] & in[74]); 
    assign layer_0[5495] = in[910] ^ in[925]; 
    assign layer_0[5496] = in[415] | in[536]; 
    assign layer_0[5497] = in[464] | in[554]; 
    assign layer_0[5498] = ~(in[328] ^ in[763]); 
    assign layer_0[5499] = ~(in[725] ^ in[296]); 
    assign layer_0[5500] = ~in[621] | (in[621] & in[619]); 
    assign layer_0[5501] = ~(in[1023] ^ in[332]); 
    assign layer_0[5502] = ~in[308]; 
    assign layer_0[5503] = in[243] ^ in[267]; 
    assign layer_0[5504] = ~in[142] | (in[142] & in[13]); 
    assign layer_0[5505] = in[855]; 
    assign layer_0[5506] = in[987] ^ in[813]; 
    assign layer_0[5507] = ~in[415]; 
    assign layer_0[5508] = in[484]; 
    assign layer_0[5509] = in[804] | in[981]; 
    assign layer_0[5510] = in[654] & ~in[983]; 
    assign layer_0[5511] = in[775] & ~in[294]; 
    assign layer_0[5512] = in[167] & in[840]; 
    assign layer_0[5513] = ~in[1014] | (in[1014] & in[763]); 
    assign layer_0[5514] = ~in[12]; 
    assign layer_0[5515] = ~in[356] | (in[783] & in[356]); 
    assign layer_0[5516] = in[441] ^ in[128]; 
    assign layer_0[5517] = in[519] | in[1018]; 
    assign layer_0[5518] = ~(in[927] | in[7]); 
    assign layer_0[5519] = in[524]; 
    assign layer_0[5520] = in[905] & in[185]; 
    assign layer_0[5521] = ~(in[585] & in[532]); 
    assign layer_0[5522] = 1'b1; 
    assign layer_0[5523] = in[901] | in[35]; 
    assign layer_0[5524] = in[868] ^ in[233]; 
    assign layer_0[5525] = ~(in[958] | in[982]); 
    assign layer_0[5526] = ~in[143]; 
    assign layer_0[5527] = ~(in[922] ^ in[967]); 
    assign layer_0[5528] = ~(in[662] ^ in[930]); 
    assign layer_0[5529] = ~(in[741] ^ in[998]); 
    assign layer_0[5530] = in[590] ^ in[207]; 
    assign layer_0[5531] = ~(in[512] & in[797]); 
    assign layer_0[5532] = ~(in[433] ^ in[452]); 
    assign layer_0[5533] = ~(in[600] ^ in[464]); 
    assign layer_0[5534] = in[905] ^ in[721]; 
    assign layer_0[5535] = ~(in[570] ^ in[656]); 
    assign layer_0[5536] = in[892] ^ in[761]; 
    assign layer_0[5537] = in[861] & ~in[889]; 
    assign layer_0[5538] = in[434] & ~in[704]; 
    assign layer_0[5539] = in[56] & ~in[588]; 
    assign layer_0[5540] = in[244] ^ in[903]; 
    assign layer_0[5541] = in[808] ^ in[3]; 
    assign layer_0[5542] = ~(in[375] ^ in[45]); 
    assign layer_0[5543] = ~in[499]; 
    assign layer_0[5544] = ~in[440]; 
    assign layer_0[5545] = in[70]; 
    assign layer_0[5546] = ~(in[500] ^ in[660]); 
    assign layer_0[5547] = ~in[580] | (in[301] & in[580]); 
    assign layer_0[5548] = in[1015] & in[483]; 
    assign layer_0[5549] = ~(in[145] ^ in[225]); 
    assign layer_0[5550] = in[628] ^ in[689]; 
    assign layer_0[5551] = ~(in[314] ^ in[952]); 
    assign layer_0[5552] = ~in[950]; 
    assign layer_0[5553] = in[858] ^ in[767]; 
    assign layer_0[5554] = ~(in[954] | in[777]); 
    assign layer_0[5555] = ~(in[987] ^ in[709]); 
    assign layer_0[5556] = in[374]; 
    assign layer_0[5557] = in[866] ^ in[744]; 
    assign layer_0[5558] = in[36] | in[31]; 
    assign layer_0[5559] = in[113] ^ in[114]; 
    assign layer_0[5560] = in[758] ^ in[759]; 
    assign layer_0[5561] = in[96] ^ in[757]; 
    assign layer_0[5562] = in[413] & ~in[276]; 
    assign layer_0[5563] = in[677] | in[578]; 
    assign layer_0[5564] = in[861] ^ in[63]; 
    assign layer_0[5565] = in[372] ^ in[253]; 
    assign layer_0[5566] = ~(in[591] ^ in[399]); 
    assign layer_0[5567] = in[632] ^ in[625]; 
    assign layer_0[5568] = ~in[868] | (in[399] & in[868]); 
    assign layer_0[5569] = in[584] | in[898]; 
    assign layer_0[5570] = in[792] & in[74]; 
    assign layer_0[5571] = in[285]; 
    assign layer_0[5572] = in[493] ^ in[355]; 
    assign layer_0[5573] = ~(in[353] & in[127]); 
    assign layer_0[5574] = ~(in[856] & in[685]); 
    assign layer_0[5575] = in[487] | in[111]; 
    assign layer_0[5576] = in[880] | in[510]; 
    assign layer_0[5577] = in[324] & ~in[682]; 
    assign layer_0[5578] = in[660] ^ in[283]; 
    assign layer_0[5579] = ~(in[850] ^ in[807]); 
    assign layer_0[5580] = in[645]; 
    assign layer_0[5581] = in[582] ^ in[306]; 
    assign layer_0[5582] = ~(in[209] ^ in[206]); 
    assign layer_0[5583] = in[587] & ~in[972]; 
    assign layer_0[5584] = in[972] & ~in[261]; 
    assign layer_0[5585] = ~(in[7] ^ in[744]); 
    assign layer_0[5586] = in[86] & ~in[946]; 
    assign layer_0[5587] = ~(in[160] ^ in[610]); 
    assign layer_0[5588] = in[748] ^ in[857]; 
    assign layer_0[5589] = ~in[687]; 
    assign layer_0[5590] = ~(in[550] ^ in[114]); 
    assign layer_0[5591] = in[445] | in[596]; 
    assign layer_0[5592] = ~in[873] | (in[873] & in[137]); 
    assign layer_0[5593] = ~(in[249] ^ in[727]); 
    assign layer_0[5594] = in[588] ^ in[886]; 
    assign layer_0[5595] = in[631] ^ in[730]; 
    assign layer_0[5596] = in[697] ^ in[253]; 
    assign layer_0[5597] = in[727] & ~in[386]; 
    assign layer_0[5598] = in[804] ^ in[283]; 
    assign layer_0[5599] = ~in[453]; 
    assign layer_0[5600] = ~(in[19] | in[735]); 
    assign layer_0[5601] = ~(in[519] | in[748]); 
    assign layer_0[5602] = ~in[698] | (in[11] & in[698]); 
    assign layer_0[5603] = in[15] & in[932]; 
    assign layer_0[5604] = ~in[424]; 
    assign layer_0[5605] = in[338] & ~in[241]; 
    assign layer_0[5606] = in[838]; 
    assign layer_0[5607] = in[965] & ~in[810]; 
    assign layer_0[5608] = ~(in[921] ^ in[920]); 
    assign layer_0[5609] = in[611] & in[450]; 
    assign layer_0[5610] = in[208] & ~in[467]; 
    assign layer_0[5611] = in[301] | in[482]; 
    assign layer_0[5612] = in[743]; 
    assign layer_0[5613] = in[884] & in[248]; 
    assign layer_0[5614] = ~(in[893] ^ in[881]); 
    assign layer_0[5615] = ~in[243] | (in[605] & in[243]); 
    assign layer_0[5616] = in[73] & ~in[163]; 
    assign layer_0[5617] = ~(in[838] ^ in[956]); 
    assign layer_0[5618] = in[41] & ~in[696]; 
    assign layer_0[5619] = ~in[411] | (in[411] & in[163]); 
    assign layer_0[5620] = ~(in[25] ^ in[822]); 
    assign layer_0[5621] = in[262] & in[204]; 
    assign layer_0[5622] = in[415] ^ in[296]; 
    assign layer_0[5623] = 1'b1; 
    assign layer_0[5624] = ~in[601] | (in[367] & in[601]); 
    assign layer_0[5625] = in[612] & ~in[871]; 
    assign layer_0[5626] = ~(in[740] ^ in[12]); 
    assign layer_0[5627] = ~in[726]; 
    assign layer_0[5628] = in[177] ^ in[443]; 
    assign layer_0[5629] = ~(in[853] & in[343]); 
    assign layer_0[5630] = in[718] & ~in[496]; 
    assign layer_0[5631] = ~in[638]; 
    assign layer_0[5632] = ~(in[821] ^ in[970]); 
    assign layer_0[5633] = ~(in[952] ^ in[156]); 
    assign layer_0[5634] = ~(in[249] ^ in[117]); 
    assign layer_0[5635] = in[617] ^ in[581]; 
    assign layer_0[5636] = ~in[92]; 
    assign layer_0[5637] = in[824] ^ in[950]; 
    assign layer_0[5638] = ~(in[420] ^ in[713]); 
    assign layer_0[5639] = ~in[888] | (in[915] & in[888]); 
    assign layer_0[5640] = ~in[760]; 
    assign layer_0[5641] = in[113]; 
    assign layer_0[5642] = in[474] & ~in[435]; 
    assign layer_0[5643] = ~(in[888] ^ in[886]); 
    assign layer_0[5644] = in[878] & in[435]; 
    assign layer_0[5645] = in[971] | in[603]; 
    assign layer_0[5646] = in[703] ^ in[400]; 
    assign layer_0[5647] = in[712] & ~in[1017]; 
    assign layer_0[5648] = ~(in[646] ^ in[474]); 
    assign layer_0[5649] = in[710] & in[900]; 
    assign layer_0[5650] = ~(in[693] ^ in[267]); 
    assign layer_0[5651] = in[691] & ~in[10]; 
    assign layer_0[5652] = ~in[57] | (in[57] & in[190]); 
    assign layer_0[5653] = in[409] & in[587]; 
    assign layer_0[5654] = in[920] | in[400]; 
    assign layer_0[5655] = ~(in[761] & in[309]); 
    assign layer_0[5656] = ~(in[1003] ^ in[259]); 
    assign layer_0[5657] = ~(in[637] & in[277]); 
    assign layer_0[5658] = ~in[206]; 
    assign layer_0[5659] = ~(in[475] ^ in[448]); 
    assign layer_0[5660] = in[808] ^ in[809]; 
    assign layer_0[5661] = in[786] ^ in[698]; 
    assign layer_0[5662] = in[12] & ~in[127]; 
    assign layer_0[5663] = in[777]; 
    assign layer_0[5664] = in[511] ^ in[370]; 
    assign layer_0[5665] = ~(in[266] ^ in[500]); 
    assign layer_0[5666] = in[596]; 
    assign layer_0[5667] = ~in[319]; 
    assign layer_0[5668] = in[902] | in[559]; 
    assign layer_0[5669] = ~in[562]; 
    assign layer_0[5670] = ~in[429] | (in[429] & in[430]); 
    assign layer_0[5671] = ~(in[581] & in[110]); 
    assign layer_0[5672] = ~in[837] | (in[837] & in[833]); 
    assign layer_0[5673] = in[692] & ~in[899]; 
    assign layer_0[5674] = ~(in[843] | in[879]); 
    assign layer_0[5675] = ~(in[671] ^ in[520]); 
    assign layer_0[5676] = ~(in[57] & in[262]); 
    assign layer_0[5677] = ~in[841] | (in[744] & in[841]); 
    assign layer_0[5678] = ~(in[807] ^ in[876]); 
    assign layer_0[5679] = ~(in[574] ^ in[968]); 
    assign layer_0[5680] = in[245] | in[720]; 
    assign layer_0[5681] = in[755] | in[208]; 
    assign layer_0[5682] = ~(in[807] ^ in[918]); 
    assign layer_0[5683] = ~(in[83] ^ in[819]); 
    assign layer_0[5684] = ~(in[666] & in[423]); 
    assign layer_0[5685] = ~(in[856] & in[215]); 
    assign layer_0[5686] = in[838] | in[274]; 
    assign layer_0[5687] = in[238] | in[759]; 
    assign layer_0[5688] = in[412] | in[683]; 
    assign layer_0[5689] = in[572] & ~in[890]; 
    assign layer_0[5690] = ~in[923]; 
    assign layer_0[5691] = ~in[680] | (in[680] & in[731]); 
    assign layer_0[5692] = in[8] & in[371]; 
    assign layer_0[5693] = in[493] ^ in[980]; 
    assign layer_0[5694] = in[759] ^ in[824]; 
    assign layer_0[5695] = in[244] & ~in[78]; 
    assign layer_0[5696] = ~in[59] | (in[59] & in[43]); 
    assign layer_0[5697] = ~in[597]; 
    assign layer_0[5698] = in[362]; 
    assign layer_0[5699] = ~in[691] | (in[899] & in[691]); 
    assign layer_0[5700] = in[185] ^ in[367]; 
    assign layer_0[5701] = ~(in[587] ^ in[875]); 
    assign layer_0[5702] = ~(in[299] & in[952]); 
    assign layer_0[5703] = in[843] ^ in[403]; 
    assign layer_0[5704] = ~in[45] | (in[45] & in[863]); 
    assign layer_0[5705] = in[939] ^ in[836]; 
    assign layer_0[5706] = ~in[496]; 
    assign layer_0[5707] = ~(in[823] | in[790]); 
    assign layer_0[5708] = ~(in[178] ^ in[623]); 
    assign layer_0[5709] = in[251] & ~in[996]; 
    assign layer_0[5710] = ~(in[222] ^ in[519]); 
    assign layer_0[5711] = ~in[7]; 
    assign layer_0[5712] = in[535] & in[715]; 
    assign layer_0[5713] = in[713] ^ in[700]; 
    assign layer_0[5714] = in[431] & ~in[643]; 
    assign layer_0[5715] = ~in[265]; 
    assign layer_0[5716] = in[379]; 
    assign layer_0[5717] = in[776] ^ in[901]; 
    assign layer_0[5718] = in[885] ^ in[4]; 
    assign layer_0[5719] = in[333]; 
    assign layer_0[5720] = in[63] & ~in[878]; 
    assign layer_0[5721] = ~in[348]; 
    assign layer_0[5722] = in[568] & ~in[483]; 
    assign layer_0[5723] = ~in[930] | (in[464] & in[930]); 
    assign layer_0[5724] = in[478] ^ in[818]; 
    assign layer_0[5725] = in[451] & in[965]; 
    assign layer_0[5726] = in[921] ^ in[730]; 
    assign layer_0[5727] = ~(in[101] ^ in[317]); 
    assign layer_0[5728] = in[711] & ~in[794]; 
    assign layer_0[5729] = ~in[555]; 
    assign layer_0[5730] = ~in[639]; 
    assign layer_0[5731] = in[985] ^ in[982]; 
    assign layer_0[5732] = ~(in[598] ^ in[518]); 
    assign layer_0[5733] = ~(in[466] ^ in[34]); 
    assign layer_0[5734] = in[855] ^ in[357]; 
    assign layer_0[5735] = in[407] & in[588]; 
    assign layer_0[5736] = in[344]; 
    assign layer_0[5737] = ~in[612] | (in[612] & in[819]); 
    assign layer_0[5738] = ~in[109]; 
    assign layer_0[5739] = ~in[336]; 
    assign layer_0[5740] = ~(in[85] & in[20]); 
    assign layer_0[5741] = ~(in[580] | in[864]); 
    assign layer_0[5742] = ~in[135]; 
    assign layer_0[5743] = ~(in[595] ^ in[253]); 
    assign layer_0[5744] = ~(in[413] & in[595]); 
    assign layer_0[5745] = 1'b0; 
    assign layer_0[5746] = in[966] ^ in[519]; 
    assign layer_0[5747] = in[159] ^ in[806]; 
    assign layer_0[5748] = ~(in[902] ^ in[431]); 
    assign layer_0[5749] = in[604]; 
    assign layer_0[5750] = ~in[692] | (in[692] & in[629]); 
    assign layer_0[5751] = in[919] & in[888]; 
    assign layer_0[5752] = in[932] ^ in[921]; 
    assign layer_0[5753] = in[708] | in[856]; 
    assign layer_0[5754] = in[677]; 
    assign layer_0[5755] = ~(in[124] ^ in[903]); 
    assign layer_0[5756] = in[63] | in[897]; 
    assign layer_0[5757] = in[678] ^ in[742]; 
    assign layer_0[5758] = in[810] ^ in[901]; 
    assign layer_0[5759] = in[911] | in[67]; 
    assign layer_0[5760] = in[299] ^ in[844]; 
    assign layer_0[5761] = in[349] & ~in[791]; 
    assign layer_0[5762] = in[912] | in[734]; 
    assign layer_0[5763] = in[94] & ~in[482]; 
    assign layer_0[5764] = ~(in[598] ^ in[615]); 
    assign layer_0[5765] = in[742] & ~in[835]; 
    assign layer_0[5766] = ~in[417] | (in[417] & in[48]); 
    assign layer_0[5767] = in[564] & ~in[351]; 
    assign layer_0[5768] = in[274] & ~in[67]; 
    assign layer_0[5769] = in[787] | in[585]; 
    assign layer_0[5770] = ~(in[855] ^ in[248]); 
    assign layer_0[5771] = in[694] & ~in[268]; 
    assign layer_0[5772] = ~(in[851] ^ in[60]); 
    assign layer_0[5773] = in[340] | in[353]; 
    assign layer_0[5774] = ~in[639]; 
    assign layer_0[5775] = ~in[319] | (in[319] & in[41]); 
    assign layer_0[5776] = ~(in[327] & in[227]); 
    assign layer_0[5777] = ~in[125] | (in[876] & in[125]); 
    assign layer_0[5778] = ~(in[945] ^ in[966]); 
    assign layer_0[5779] = ~in[701] | (in[3] & in[701]); 
    assign layer_0[5780] = ~(in[957] | in[433]); 
    assign layer_0[5781] = ~in[594]; 
    assign layer_0[5782] = ~(in[227] ^ in[204]); 
    assign layer_0[5783] = ~(in[315] | in[263]); 
    assign layer_0[5784] = in[847] | in[759]; 
    assign layer_0[5785] = in[262] | in[867]; 
    assign layer_0[5786] = ~(in[477] ^ in[954]); 
    assign layer_0[5787] = in[2] & ~in[493]; 
    assign layer_0[5788] = in[161] | in[518]; 
    assign layer_0[5789] = ~(in[899] ^ in[997]); 
    assign layer_0[5790] = ~(in[657] & in[616]); 
    assign layer_0[5791] = ~(in[475] & in[820]); 
    assign layer_0[5792] = in[443] ^ in[663]; 
    assign layer_0[5793] = in[612] ^ in[603]; 
    assign layer_0[5794] = in[437] & ~in[488]; 
    assign layer_0[5795] = ~(in[917] ^ in[762]); 
    assign layer_0[5796] = in[290] ^ in[266]; 
    assign layer_0[5797] = in[885] | in[339]; 
    assign layer_0[5798] = in[523] | in[516]; 
    assign layer_0[5799] = ~(in[4] ^ in[504]); 
    assign layer_0[5800] = in[583] & ~in[851]; 
    assign layer_0[5801] = in[132] & ~in[572]; 
    assign layer_0[5802] = in[1018] | in[386]; 
    assign layer_0[5803] = ~in[176] | (in[176] & in[257]); 
    assign layer_0[5804] = ~in[858]; 
    assign layer_0[5805] = ~in[423] | (in[423] & in[45]); 
    assign layer_0[5806] = in[624]; 
    assign layer_0[5807] = in[162] & in[762]; 
    assign layer_0[5808] = in[97] ^ in[392]; 
    assign layer_0[5809] = ~(in[968] ^ in[276]); 
    assign layer_0[5810] = ~in[100] | (in[100] & in[912]); 
    assign layer_0[5811] = ~in[169] | (in[318] & in[169]); 
    assign layer_0[5812] = in[173] | in[496]; 
    assign layer_0[5813] = ~in[159] | (in[159] & in[476]); 
    assign layer_0[5814] = ~(in[327] ^ in[676]); 
    assign layer_0[5815] = in[569]; 
    assign layer_0[5816] = ~in[720]; 
    assign layer_0[5817] = in[493] ^ in[302]; 
    assign layer_0[5818] = ~(in[607] | in[757]); 
    assign layer_0[5819] = ~in[956]; 
    assign layer_0[5820] = ~in[808] | (in[808] & in[821]); 
    assign layer_0[5821] = ~in[851]; 
    assign layer_0[5822] = ~(in[823] ^ in[127]); 
    assign layer_0[5823] = in[998] & ~in[884]; 
    assign layer_0[5824] = ~(in[6] ^ in[176]); 
    assign layer_0[5825] = ~(in[179] ^ in[720]); 
    assign layer_0[5826] = in[466] | in[467]; 
    assign layer_0[5827] = in[589]; 
    assign layer_0[5828] = in[102] | in[890]; 
    assign layer_0[5829] = ~(in[175] | in[844]); 
    assign layer_0[5830] = ~(in[264] ^ in[555]); 
    assign layer_0[5831] = in[467] ^ in[676]; 
    assign layer_0[5832] = in[424]; 
    assign layer_0[5833] = ~(in[120] & in[476]); 
    assign layer_0[5834] = ~in[316] | (in[316] & in[111]); 
    assign layer_0[5835] = in[210] ^ in[615]; 
    assign layer_0[5836] = ~in[758] | (in[758] & in[259]); 
    assign layer_0[5837] = ~(in[146] ^ in[776]); 
    assign layer_0[5838] = in[420] ^ in[341]; 
    assign layer_0[5839] = in[167] & ~in[920]; 
    assign layer_0[5840] = in[1000] | in[557]; 
    assign layer_0[5841] = ~(in[17] ^ in[1000]); 
    assign layer_0[5842] = ~in[886]; 
    assign layer_0[5843] = in[935] & ~in[824]; 
    assign layer_0[5844] = in[899] & ~in[262]; 
    assign layer_0[5845] = ~(in[536] | in[44]); 
    assign layer_0[5846] = ~(in[459] ^ in[794]); 
    assign layer_0[5847] = in[310] & ~in[189]; 
    assign layer_0[5848] = in[793]; 
    assign layer_0[5849] = in[754] | in[201]; 
    assign layer_0[5850] = in[844]; 
    assign layer_0[5851] = in[551] & ~in[63]; 
    assign layer_0[5852] = ~(in[955] ^ in[685]); 
    assign layer_0[5853] = in[856] ^ in[937]; 
    assign layer_0[5854] = in[856] | in[236]; 
    assign layer_0[5855] = ~(in[836] ^ in[772]); 
    assign layer_0[5856] = ~(in[220] ^ in[571]); 
    assign layer_0[5857] = ~in[373] | (in[264] & in[373]); 
    assign layer_0[5858] = 1'b0; 
    assign layer_0[5859] = in[85] | in[596]; 
    assign layer_0[5860] = in[602] ^ in[966]; 
    assign layer_0[5861] = ~(in[427] ^ in[336]); 
    assign layer_0[5862] = ~(in[602] ^ in[138]); 
    assign layer_0[5863] = ~(in[839] ^ in[380]); 
    assign layer_0[5864] = in[268]; 
    assign layer_0[5865] = ~(in[792] ^ in[953]); 
    assign layer_0[5866] = in[519] ^ in[548]; 
    assign layer_0[5867] = in[144] ^ in[450]; 
    assign layer_0[5868] = ~(in[218] & in[682]); 
    assign layer_0[5869] = ~(in[954] ^ in[241]); 
    assign layer_0[5870] = ~in[922] | (in[10] & in[922]); 
    assign layer_0[5871] = ~in[262]; 
    assign layer_0[5872] = ~(in[857] ^ in[260]); 
    assign layer_0[5873] = in[565]; 
    assign layer_0[5874] = in[307] ^ in[517]; 
    assign layer_0[5875] = in[563] ^ in[486]; 
    assign layer_0[5876] = ~(in[489] & in[490]); 
    assign layer_0[5877] = ~(in[749] ^ in[838]); 
    assign layer_0[5878] = in[496]; 
    assign layer_0[5879] = ~(in[704] | in[285]); 
    assign layer_0[5880] = ~(in[950] ^ in[933]); 
    assign layer_0[5881] = ~(in[324] | in[915]); 
    assign layer_0[5882] = in[729] ^ in[967]; 
    assign layer_0[5883] = ~in[310] | (in[310] & in[79]); 
    assign layer_0[5884] = in[974] ^ in[714]; 
    assign layer_0[5885] = in[327] ^ in[607]; 
    assign layer_0[5886] = ~(in[524] ^ in[557]); 
    assign layer_0[5887] = in[674] ^ in[534]; 
    assign layer_0[5888] = ~(in[278] ^ in[667]); 
    assign layer_0[5889] = in[536] ^ in[533]; 
    assign layer_0[5890] = ~in[40] | (in[40] & in[517]); 
    assign layer_0[5891] = in[461] ^ in[237]; 
    assign layer_0[5892] = in[591] ^ in[296]; 
    assign layer_0[5893] = ~(in[875] ^ in[921]); 
    assign layer_0[5894] = ~(in[65] | in[111]); 
    assign layer_0[5895] = ~(in[717] | in[850]); 
    assign layer_0[5896] = ~(in[619] ^ in[1015]); 
    assign layer_0[5897] = ~(in[608] | in[938]); 
    assign layer_0[5898] = in[862] ^ in[218]; 
    assign layer_0[5899] = ~in[648]; 
    assign layer_0[5900] = ~in[300]; 
    assign layer_0[5901] = in[886] ^ in[923]; 
    assign layer_0[5902] = in[725]; 
    assign layer_0[5903] = ~(in[430] ^ in[884]); 
    assign layer_0[5904] = ~(in[910] ^ in[448]); 
    assign layer_0[5905] = in[805]; 
    assign layer_0[5906] = in[181]; 
    assign layer_0[5907] = ~in[364] | (in[364] & in[262]); 
    assign layer_0[5908] = ~(in[435] ^ in[157]); 
    assign layer_0[5909] = ~in[761] | (in[51] & in[761]); 
    assign layer_0[5910] = in[150]; 
    assign layer_0[5911] = ~in[878] | (in[911] & in[878]); 
    assign layer_0[5912] = in[8] & ~in[545]; 
    assign layer_0[5913] = in[6] | in[834]; 
    assign layer_0[5914] = in[12] & ~in[939]; 
    assign layer_0[5915] = ~(in[313] & in[999]); 
    assign layer_0[5916] = in[698]; 
    assign layer_0[5917] = ~(in[687] | in[680]); 
    assign layer_0[5918] = ~(in[950] & in[668]); 
    assign layer_0[5919] = in[823]; 
    assign layer_0[5920] = in[760] & ~in[333]; 
    assign layer_0[5921] = in[534] ^ in[822]; 
    assign layer_0[5922] = in[947] & ~in[245]; 
    assign layer_0[5923] = ~(in[1000] ^ in[984]); 
    assign layer_0[5924] = ~(in[353] ^ in[491]); 
    assign layer_0[5925] = in[318] ^ in[626]; 
    assign layer_0[5926] = ~(in[715] ^ in[436]); 
    assign layer_0[5927] = ~(in[565] ^ in[548]); 
    assign layer_0[5928] = ~(in[277] ^ in[490]); 
    assign layer_0[5929] = ~(in[915] | in[194]); 
    assign layer_0[5930] = 1'b0; 
    assign layer_0[5931] = ~(in[868] & in[966]); 
    assign layer_0[5932] = in[537] & in[877]; 
    assign layer_0[5933] = in[132] ^ in[857]; 
    assign layer_0[5934] = in[590] ^ in[893]; 
    assign layer_0[5935] = ~(in[474] | in[578]); 
    assign layer_0[5936] = in[259] & in[323]; 
    assign layer_0[5937] = in[538] | in[360]; 
    assign layer_0[5938] = in[984] ^ in[947]; 
    assign layer_0[5939] = in[567] & in[597]; 
    assign layer_0[5940] = ~(in[503] ^ in[748]); 
    assign layer_0[5941] = in[371] ^ in[407]; 
    assign layer_0[5942] = ~(in[89] & in[762]); 
    assign layer_0[5943] = ~(in[10] ^ in[935]); 
    assign layer_0[5944] = in[332] ^ in[982]; 
    assign layer_0[5945] = ~in[45] | (in[947] & in[45]); 
    assign layer_0[5946] = in[775]; 
    assign layer_0[5947] = ~(in[869] ^ in[842]); 
    assign layer_0[5948] = in[966] & ~in[512]; 
    assign layer_0[5949] = in[794] & ~in[17]; 
    assign layer_0[5950] = ~in[341]; 
    assign layer_0[5951] = in[293] ^ in[954]; 
    assign layer_0[5952] = in[583] & in[191]; 
    assign layer_0[5953] = ~(in[483] ^ in[730]); 
    assign layer_0[5954] = ~in[829]; 
    assign layer_0[5955] = in[150]; 
    assign layer_0[5956] = in[583] & ~in[945]; 
    assign layer_0[5957] = in[370]; 
    assign layer_0[5958] = in[587] & in[572]; 
    assign layer_0[5959] = ~in[360] | (in[893] & in[360]); 
    assign layer_0[5960] = in[849] | in[63]; 
    assign layer_0[5961] = 1'b1; 
    assign layer_0[5962] = ~in[428] | (in[428] & in[870]); 
    assign layer_0[5963] = in[425] ^ in[3]; 
    assign layer_0[5964] = ~in[605]; 
    assign layer_0[5965] = in[536] ^ in[731]; 
    assign layer_0[5966] = ~in[903]; 
    assign layer_0[5967] = in[218] & ~in[557]; 
    assign layer_0[5968] = in[429] & ~in[291]; 
    assign layer_0[5969] = in[554] & ~in[653]; 
    assign layer_0[5970] = in[898] & ~in[225]; 
    assign layer_0[5971] = ~(in[70] | in[704]); 
    assign layer_0[5972] = in[680]; 
    assign layer_0[5973] = in[330] ^ in[717]; 
    assign layer_0[5974] = in[376] & ~in[712]; 
    assign layer_0[5975] = ~(in[810] ^ in[243]); 
    assign layer_0[5976] = ~(in[334] | in[334]); 
    assign layer_0[5977] = in[193] ^ in[775]; 
    assign layer_0[5978] = in[762] ^ in[886]; 
    assign layer_0[5979] = in[357] | in[86]; 
    assign layer_0[5980] = ~(in[299] ^ in[952]); 
    assign layer_0[5981] = in[226]; 
    assign layer_0[5982] = in[526] | in[603]; 
    assign layer_0[5983] = ~in[979]; 
    assign layer_0[5984] = in[462] & ~in[713]; 
    assign layer_0[5985] = in[308] ^ in[678]; 
    assign layer_0[5986] = ~(in[418] ^ in[226]); 
    assign layer_0[5987] = in[641] & ~in[576]; 
    assign layer_0[5988] = ~(in[538] ^ in[555]); 
    assign layer_0[5989] = in[10] ^ in[296]; 
    assign layer_0[5990] = ~(in[731] ^ in[275]); 
    assign layer_0[5991] = ~(in[857] ^ in[356]); 
    assign layer_0[5992] = in[308] | in[279]; 
    assign layer_0[5993] = ~(in[289] | in[284]); 
    assign layer_0[5994] = ~in[938] | (in[938] & in[25]); 
    assign layer_0[5995] = ~(in[591] | in[988]); 
    assign layer_0[5996] = ~in[808] | (in[5] & in[808]); 
    assign layer_0[5997] = ~(in[882] ^ in[888]); 
    assign layer_0[5998] = ~(in[692] ^ in[94]); 
    assign layer_0[5999] = ~(in[445] & in[36]); 
    assign layer_0[6000] = in[889] ^ in[158]; 
    assign layer_0[6001] = in[50] & in[732]; 
    assign layer_0[6002] = in[227] & ~in[651]; 
    assign layer_0[6003] = ~in[619] | (in[839] & in[619]); 
    assign layer_0[6004] = ~(in[431] ^ in[593]); 
    assign layer_0[6005] = in[302] & in[829]; 
    assign layer_0[6006] = in[853]; 
    assign layer_0[6007] = in[46] & in[198]; 
    assign layer_0[6008] = in[632] & in[1018]; 
    assign layer_0[6009] = ~(in[285] ^ in[746]); 
    assign layer_0[6010] = in[122]; 
    assign layer_0[6011] = ~(in[453] ^ in[927]); 
    assign layer_0[6012] = in[35] ^ in[704]; 
    assign layer_0[6013] = ~(in[604] | in[577]); 
    assign layer_0[6014] = in[928] & ~in[501]; 
    assign layer_0[6015] = in[356] & ~in[601]; 
    assign layer_0[6016] = ~(in[439] ^ in[230]); 
    assign layer_0[6017] = ~(in[555] ^ in[1001]); 
    assign layer_0[6018] = ~in[521] | (in[688] & in[521]); 
    assign layer_0[6019] = in[424] ^ in[683]; 
    assign layer_0[6020] = ~in[288] | (in[288] & in[433]); 
    assign layer_0[6021] = in[883]; 
    assign layer_0[6022] = in[520] & ~in[888]; 
    assign layer_0[6023] = ~in[56] | (in[1003] & in[56]); 
    assign layer_0[6024] = ~(in[520] | in[921]); 
    assign layer_0[6025] = in[640] & ~in[282]; 
    assign layer_0[6026] = ~in[905] | (in[722] & in[905]); 
    assign layer_0[6027] = ~(in[76] | in[357]); 
    assign layer_0[6028] = ~in[875] | (in[342] & in[875]); 
    assign layer_0[6029] = in[580] ^ in[99]; 
    assign layer_0[6030] = in[902] ^ in[983]; 
    assign layer_0[6031] = ~(in[936] ^ in[950]); 
    assign layer_0[6032] = in[464] | in[556]; 
    assign layer_0[6033] = in[915] & ~in[499]; 
    assign layer_0[6034] = ~(in[707] ^ in[459]); 
    assign layer_0[6035] = in[930] | in[554]; 
    assign layer_0[6036] = ~(in[924] ^ in[724]); 
    assign layer_0[6037] = ~in[1015]; 
    assign layer_0[6038] = ~in[818] | (in[890] & in[818]); 
    assign layer_0[6039] = ~(in[745] ^ in[502]); 
    assign layer_0[6040] = ~in[271] | (in[271] & in[418]); 
    assign layer_0[6041] = ~(in[926] ^ in[940]); 
    assign layer_0[6042] = ~(in[665] & in[617]); 
    assign layer_0[6043] = ~(in[897] | in[369]); 
    assign layer_0[6044] = in[1000]; 
    assign layer_0[6045] = in[424] & in[396]; 
    assign layer_0[6046] = ~(in[587] ^ in[722]); 
    assign layer_0[6047] = in[410] & ~in[793]; 
    assign layer_0[6048] = ~(in[987] | in[737]); 
    assign layer_0[6049] = in[196] & ~in[716]; 
    assign layer_0[6050] = in[471] ^ in[916]; 
    assign layer_0[6051] = in[936] ^ in[507]; 
    assign layer_0[6052] = ~(in[810] ^ in[582]); 
    assign layer_0[6053] = in[7]; 
    assign layer_0[6054] = in[983]; 
    assign layer_0[6055] = ~(in[826] | in[915]); 
    assign layer_0[6056] = in[341] & ~in[33]; 
    assign layer_0[6057] = 1'b1; 
    assign layer_0[6058] = in[842] | in[438]; 
    assign layer_0[6059] = ~(in[795] | in[963]); 
    assign layer_0[6060] = in[397] & in[483]; 
    assign layer_0[6061] = in[855]; 
    assign layer_0[6062] = in[3] & ~in[831]; 
    assign layer_0[6063] = in[1018] ^ in[854]; 
    assign layer_0[6064] = in[119] ^ in[229]; 
    assign layer_0[6065] = ~(in[852] | in[581]); 
    assign layer_0[6066] = in[638] ^ in[451]; 
    assign layer_0[6067] = ~(in[463] | in[825]); 
    assign layer_0[6068] = in[748] | in[290]; 
    assign layer_0[6069] = ~in[333] | (in[762] & in[333]); 
    assign layer_0[6070] = ~in[997] | (in[997] & in[4]); 
    assign layer_0[6071] = in[891] & ~in[221]; 
    assign layer_0[6072] = in[1] & in[437]; 
    assign layer_0[6073] = ~in[419]; 
    assign layer_0[6074] = in[483] ^ in[594]; 
    assign layer_0[6075] = ~(in[413] & in[696]); 
    assign layer_0[6076] = in[483] & in[966]; 
    assign layer_0[6077] = ~(in[432] & in[145]); 
    assign layer_0[6078] = 1'b0; 
    assign layer_0[6079] = ~(in[131] ^ in[806]); 
    assign layer_0[6080] = ~(in[857] | in[417]); 
    assign layer_0[6081] = in[262] & ~in[962]; 
    assign layer_0[6082] = ~(in[466] | in[1001]); 
    assign layer_0[6083] = ~in[963] | (in[963] & in[954]); 
    assign layer_0[6084] = in[743] & in[599]; 
    assign layer_0[6085] = in[250]; 
    assign layer_0[6086] = ~(in[362] & in[174]); 
    assign layer_0[6087] = ~(in[77] & in[601]); 
    assign layer_0[6088] = ~in[731]; 
    assign layer_0[6089] = ~in[747] | (in[747] & in[92]); 
    assign layer_0[6090] = in[949]; 
    assign layer_0[6091] = in[669] ^ in[231]; 
    assign layer_0[6092] = ~in[474] | (in[474] & in[262]); 
    assign layer_0[6093] = in[283]; 
    assign layer_0[6094] = ~(in[354] & in[875]); 
    assign layer_0[6095] = 1'b0; 
    assign layer_0[6096] = ~in[8] | (in[630] & in[8]); 
    assign layer_0[6097] = in[415] | in[771]; 
    assign layer_0[6098] = in[885] ^ in[350]; 
    assign layer_0[6099] = in[621] ^ in[142]; 
    assign layer_0[6100] = ~(in[306] ^ in[482]); 
    assign layer_0[6101] = in[971] ^ in[840]; 
    assign layer_0[6102] = ~in[665] | (in[445] & in[665]); 
    assign layer_0[6103] = ~(in[83] ^ in[979]); 
    assign layer_0[6104] = in[776] ^ in[938]; 
    assign layer_0[6105] = in[312] & ~in[464]; 
    assign layer_0[6106] = ~in[96]; 
    assign layer_0[6107] = in[761] ^ in[28]; 
    assign layer_0[6108] = ~(in[386] ^ in[243]); 
    assign layer_0[6109] = ~(in[607] ^ in[313]); 
    assign layer_0[6110] = in[266] & in[40]; 
    assign layer_0[6111] = in[62] | in[1003]; 
    assign layer_0[6112] = in[366]; 
    assign layer_0[6113] = ~(in[906] ^ in[683]); 
    assign layer_0[6114] = ~in[796]; 
    assign layer_0[6115] = in[965] ^ in[413]; 
    assign layer_0[6116] = ~in[573] | (in[334] & in[573]); 
    assign layer_0[6117] = in[569] ^ in[601]; 
    assign layer_0[6118] = in[535] ^ in[787]; 
    assign layer_0[6119] = in[548] ^ in[853]; 
    assign layer_0[6120] = ~(in[111] | in[520]); 
    assign layer_0[6121] = in[317]; 
    assign layer_0[6122] = in[910] & ~in[725]; 
    assign layer_0[6123] = ~(in[484] ^ in[950]); 
    assign layer_0[6124] = ~in[947]; 
    assign layer_0[6125] = ~(in[628] | in[723]); 
    assign layer_0[6126] = ~(in[543] ^ in[213]); 
    assign layer_0[6127] = in[632] ^ in[281]; 
    assign layer_0[6128] = in[696] & ~in[982]; 
    assign layer_0[6129] = ~in[55]; 
    assign layer_0[6130] = 1'b1; 
    assign layer_0[6131] = ~(in[415] ^ in[144]); 
    assign layer_0[6132] = ~(in[484] | in[932]); 
    assign layer_0[6133] = ~in[810] | (in[810] & in[949]); 
    assign layer_0[6134] = in[918] | in[742]; 
    assign layer_0[6135] = ~in[675]; 
    assign layer_0[6136] = ~in[345] | (in[351] & in[345]); 
    assign layer_0[6137] = in[467] ^ in[874]; 
    assign layer_0[6138] = in[190] | in[889]; 
    assign layer_0[6139] = in[634] & ~in[589]; 
    assign layer_0[6140] = in[681] & ~in[276]; 
    assign layer_0[6141] = in[901] | in[542]; 
    assign layer_0[6142] = in[892]; 
    assign layer_0[6143] = ~(in[116] & in[144]); 
    assign layer_0[6144] = in[300] ^ in[533]; 
    assign layer_0[6145] = in[973] ^ in[724]; 
    assign layer_0[6146] = in[952] ^ in[259]; 
    assign layer_0[6147] = ~in[294] | (in[1014] & in[294]); 
    assign layer_0[6148] = in[709] & in[535]; 
    assign layer_0[6149] = in[986] ^ in[200]; 
    assign layer_0[6150] = ~in[940] | (in[864] & in[940]); 
    assign layer_0[6151] = ~in[777]; 
    assign layer_0[6152] = ~in[616]; 
    assign layer_0[6153] = in[835] | in[729]; 
    assign layer_0[6154] = in[457] & ~in[984]; 
    assign layer_0[6155] = in[859] ^ in[50]; 
    assign layer_0[6156] = ~(in[0] ^ in[739]); 
    assign layer_0[6157] = in[842] & ~in[341]; 
    assign layer_0[6158] = in[261] ^ in[507]; 
    assign layer_0[6159] = in[24] & in[177]; 
    assign layer_0[6160] = in[616]; 
    assign layer_0[6161] = in[260] ^ in[500]; 
    assign layer_0[6162] = in[369] & ~in[855]; 
    assign layer_0[6163] = ~(in[365] ^ in[853]); 
    assign layer_0[6164] = ~(in[938] ^ in[122]); 
    assign layer_0[6165] = ~in[718]; 
    assign layer_0[6166] = in[870] & in[401]; 
    assign layer_0[6167] = ~(in[761] ^ in[356]); 
    assign layer_0[6168] = in[82]; 
    assign layer_0[6169] = in[969] ^ in[633]; 
    assign layer_0[6170] = ~(in[915] ^ in[669]); 
    assign layer_0[6171] = ~in[903] | (in[844] & in[903]); 
    assign layer_0[6172] = ~(in[805] ^ in[762]); 
    assign layer_0[6173] = ~(in[460] & in[908]); 
    assign layer_0[6174] = in[699] & in[114]; 
    assign layer_0[6175] = in[40] & ~in[993]; 
    assign layer_0[6176] = ~in[951]; 
    assign layer_0[6177] = 1'b0; 
    assign layer_0[6178] = ~(in[677] ^ in[726]); 
    assign layer_0[6179] = in[485] ^ in[35]; 
    assign layer_0[6180] = in[612] & ~in[446]; 
    assign layer_0[6181] = 1'b0; 
    assign layer_0[6182] = 1'b0; 
    assign layer_0[6183] = in[235] & ~in[969]; 
    assign layer_0[6184] = ~in[910] | (in[773] & in[910]); 
    assign layer_0[6185] = in[840] ^ in[999]; 
    assign layer_0[6186] = ~(in[187] & in[572]); 
    assign layer_0[6187] = ~(in[266] & in[231]); 
    assign layer_0[6188] = in[253] ^ in[411]; 
    assign layer_0[6189] = in[716] ^ in[684]; 
    assign layer_0[6190] = in[850] | in[61]; 
    assign layer_0[6191] = in[76] & ~in[961]; 
    assign layer_0[6192] = ~in[934]; 
    assign layer_0[6193] = ~(in[15] | in[113]); 
    assign layer_0[6194] = in[614] & ~in[825]; 
    assign layer_0[6195] = in[517]; 
    assign layer_0[6196] = in[847] & ~in[701]; 
    assign layer_0[6197] = in[618] ^ in[650]; 
    assign layer_0[6198] = ~(in[477] ^ in[51]); 
    assign layer_0[6199] = in[19] & ~in[584]; 
    assign layer_0[6200] = in[142]; 
    assign layer_0[6201] = ~(in[460] | in[129]); 
    assign layer_0[6202] = in[646] ^ in[451]; 
    assign layer_0[6203] = in[132] | in[321]; 
    assign layer_0[6204] = in[243] & in[323]; 
    assign layer_0[6205] = in[233] ^ in[79]; 
    assign layer_0[6206] = ~(in[724] ^ in[420]); 
    assign layer_0[6207] = ~(in[198] ^ in[218]); 
    assign layer_0[6208] = in[28] & in[357]; 
    assign layer_0[6209] = in[935] & ~in[3]; 
    assign layer_0[6210] = ~in[966] | (in[850] & in[966]); 
    assign layer_0[6211] = in[840]; 
    assign layer_0[6212] = ~in[485] | (in[811] & in[485]); 
    assign layer_0[6213] = in[633]; 
    assign layer_0[6214] = ~(in[69] ^ in[897]); 
    assign layer_0[6215] = ~(in[227] ^ in[193]); 
    assign layer_0[6216] = in[725] ^ in[995]; 
    assign layer_0[6217] = ~(in[534] ^ in[795]); 
    assign layer_0[6218] = ~(in[888] ^ in[984]); 
    assign layer_0[6219] = ~in[1001]; 
    assign layer_0[6220] = ~(in[268] ^ in[44]); 
    assign layer_0[6221] = in[587] ^ in[612]; 
    assign layer_0[6222] = ~in[948]; 
    assign layer_0[6223] = in[617]; 
    assign layer_0[6224] = ~(in[749] ^ in[662]); 
    assign layer_0[6225] = in[21] ^ in[294]; 
    assign layer_0[6226] = ~in[500] | (in[500] & in[902]); 
    assign layer_0[6227] = in[901] ^ in[448]; 
    assign layer_0[6228] = in[285]; 
    assign layer_0[6229] = in[749] ^ in[647]; 
    assign layer_0[6230] = in[467] ^ in[650]; 
    assign layer_0[6231] = 1'b0; 
    assign layer_0[6232] = in[338]; 
    assign layer_0[6233] = in[231]; 
    assign layer_0[6234] = in[406] & ~in[628]; 
    assign layer_0[6235] = ~in[744]; 
    assign layer_0[6236] = in[932] | in[810]; 
    assign layer_0[6237] = ~in[32] | (in[32] & in[971]); 
    assign layer_0[6238] = ~(in[32] & in[23]); 
    assign layer_0[6239] = in[612] ^ in[28]; 
    assign layer_0[6240] = ~in[99]; 
    assign layer_0[6241] = in[489]; 
    assign layer_0[6242] = in[268] & ~in[15]; 
    assign layer_0[6243] = in[745]; 
    assign layer_0[6244] = in[951] ^ in[969]; 
    assign layer_0[6245] = ~(in[744] ^ in[742]); 
    assign layer_0[6246] = in[328] ^ in[200]; 
    assign layer_0[6247] = ~(in[916] ^ in[984]); 
    assign layer_0[6248] = ~(in[911] | in[448]); 
    assign layer_0[6249] = in[502] ^ in[336]; 
    assign layer_0[6250] = ~(in[809] & in[410]); 
    assign layer_0[6251] = ~in[404] | (in[157] & in[404]); 
    assign layer_0[6252] = ~in[386]; 
    assign layer_0[6253] = ~(in[891] | in[689]); 
    assign layer_0[6254] = ~(in[872] ^ in[887]); 
    assign layer_0[6255] = ~in[655]; 
    assign layer_0[6256] = ~in[174] | (in[174] & in[208]); 
    assign layer_0[6257] = in[373] ^ in[54]; 
    assign layer_0[6258] = ~(in[860] ^ in[772]); 
    assign layer_0[6259] = in[431] ^ in[534]; 
    assign layer_0[6260] = in[109] | in[1018]; 
    assign layer_0[6261] = in[964] & ~in[942]; 
    assign layer_0[6262] = in[307]; 
    assign layer_0[6263] = ~in[963] | (in[963] & in[1019]); 
    assign layer_0[6264] = in[126] ^ in[956]; 
    assign layer_0[6265] = ~(in[325] ^ in[921]); 
    assign layer_0[6266] = in[662]; 
    assign layer_0[6267] = in[921] | in[752]; 
    assign layer_0[6268] = in[860] & ~in[972]; 
    assign layer_0[6269] = ~in[873] | (in[873] & in[879]); 
    assign layer_0[6270] = in[498] | in[991]; 
    assign layer_0[6271] = in[221]; 
    assign layer_0[6272] = in[621] ^ in[604]; 
    assign layer_0[6273] = ~in[43] | (in[376] & in[43]); 
    assign layer_0[6274] = in[838] ^ in[837]; 
    assign layer_0[6275] = in[449] & ~in[99]; 
    assign layer_0[6276] = ~(in[917] & in[676]); 
    assign layer_0[6277] = in[985] ^ in[868]; 
    assign layer_0[6278] = ~(in[602] & in[597]); 
    assign layer_0[6279] = ~(in[540] ^ in[126]); 
    assign layer_0[6280] = ~(in[854] ^ in[967]); 
    assign layer_0[6281] = in[275]; 
    assign layer_0[6282] = ~in[100] | (in[100] & in[947]); 
    assign layer_0[6283] = ~(in[430] ^ in[570]); 
    assign layer_0[6284] = ~in[11] | (in[643] & in[11]); 
    assign layer_0[6285] = in[262] & ~in[12]; 
    assign layer_0[6286] = ~in[212]; 
    assign layer_0[6287] = ~(in[476] ^ in[901]); 
    assign layer_0[6288] = ~(in[12] ^ in[332]); 
    assign layer_0[6289] = in[583] | in[203]; 
    assign layer_0[6290] = ~(in[388] ^ in[375]); 
    assign layer_0[6291] = in[64] | in[517]; 
    assign layer_0[6292] = in[682] ^ in[603]; 
    assign layer_0[6293] = in[22]; 
    assign layer_0[6294] = ~(in[299] ^ in[520]); 
    assign layer_0[6295] = ~(in[743] ^ in[117]); 
    assign layer_0[6296] = 1'b1; 
    assign layer_0[6297] = ~(in[753] | in[599]); 
    assign layer_0[6298] = in[154] & ~in[91]; 
    assign layer_0[6299] = ~(in[681] | in[941]); 
    assign layer_0[6300] = in[932]; 
    assign layer_0[6301] = in[581] ^ in[936]; 
    assign layer_0[6302] = ~in[663]; 
    assign layer_0[6303] = ~(in[963] ^ in[692]); 
    assign layer_0[6304] = in[482] | in[318]; 
    assign layer_0[6305] = in[919] ^ in[226]; 
    assign layer_0[6306] = in[631] | in[7]; 
    assign layer_0[6307] = in[25]; 
    assign layer_0[6308] = ~in[378] | (in[914] & in[378]); 
    assign layer_0[6309] = in[911] ^ in[589]; 
    assign layer_0[6310] = in[392]; 
    assign layer_0[6311] = in[604] & ~in[714]; 
    assign layer_0[6312] = in[715] | in[585]; 
    assign layer_0[6313] = ~(in[809] | in[477]); 
    assign layer_0[6314] = in[220] & ~in[444]; 
    assign layer_0[6315] = ~(in[576] | in[725]); 
    assign layer_0[6316] = ~in[311]; 
    assign layer_0[6317] = in[276] ^ in[12]; 
    assign layer_0[6318] = ~(in[61] ^ in[329]); 
    assign layer_0[6319] = ~in[812] | (in[812] & in[964]); 
    assign layer_0[6320] = in[851] & ~in[550]; 
    assign layer_0[6321] = in[442] | in[158]; 
    assign layer_0[6322] = in[451]; 
    assign layer_0[6323] = in[377] & ~in[368]; 
    assign layer_0[6324] = ~(in[461] ^ in[823]); 
    assign layer_0[6325] = in[234] ^ in[174]; 
    assign layer_0[6326] = in[215] ^ in[660]; 
    assign layer_0[6327] = in[113] & ~in[133]; 
    assign layer_0[6328] = ~(in[450] & in[745]); 
    assign layer_0[6329] = in[893] ^ in[966]; 
    assign layer_0[6330] = in[71] ^ in[860]; 
    assign layer_0[6331] = ~(in[984] & in[564]); 
    assign layer_0[6332] = ~(in[337] & in[101]); 
    assign layer_0[6333] = 1'b0; 
    assign layer_0[6334] = in[459] ^ in[901]; 
    assign layer_0[6335] = ~in[323]; 
    assign layer_0[6336] = in[599] | in[319]; 
    assign layer_0[6337] = in[534] ^ in[913]; 
    assign layer_0[6338] = ~(in[536] ^ in[807]); 
    assign layer_0[6339] = in[157]; 
    assign layer_0[6340] = ~in[856] | (in[856] & in[824]); 
    assign layer_0[6341] = ~(in[639] ^ in[194]); 
    assign layer_0[6342] = in[669] ^ in[1004]; 
    assign layer_0[6343] = in[818] | in[716]; 
    assign layer_0[6344] = ~(in[63] ^ in[732]); 
    assign layer_0[6345] = ~(in[520] & in[565]); 
    assign layer_0[6346] = in[422] ^ in[16]; 
    assign layer_0[6347] = in[837] & ~in[317]; 
    assign layer_0[6348] = ~(in[858] ^ in[1015]); 
    assign layer_0[6349] = in[45] & ~in[848]; 
    assign layer_0[6350] = ~(in[152] ^ in[15]); 
    assign layer_0[6351] = in[247] & in[521]; 
    assign layer_0[6352] = in[900] & ~in[707]; 
    assign layer_0[6353] = in[726] ^ in[534]; 
    assign layer_0[6354] = ~(in[282] | in[776]); 
    assign layer_0[6355] = in[821] ^ in[174]; 
    assign layer_0[6356] = in[941] ^ in[568]; 
    assign layer_0[6357] = in[519] & ~in[260]; 
    assign layer_0[6358] = ~(in[947] ^ in[840]); 
    assign layer_0[6359] = in[854] & in[635]; 
    assign layer_0[6360] = in[696] ^ in[373]; 
    assign layer_0[6361] = ~(in[742] ^ in[741]); 
    assign layer_0[6362] = ~in[747] | (in[917] & in[747]); 
    assign layer_0[6363] = ~(in[896] ^ in[332]); 
    assign layer_0[6364] = in[838] & ~in[903]; 
    assign layer_0[6365] = ~(in[280] | in[437]); 
    assign layer_0[6366] = in[1000] ^ in[952]; 
    assign layer_0[6367] = ~(in[257] & in[286]); 
    assign layer_0[6368] = in[298] | in[626]; 
    assign layer_0[6369] = ~in[659] | (in[659] & in[129]); 
    assign layer_0[6370] = in[201] & in[997]; 
    assign layer_0[6371] = in[270] ^ in[396]; 
    assign layer_0[6372] = in[839] ^ in[840]; 
    assign layer_0[6373] = in[602] & ~in[968]; 
    assign layer_0[6374] = in[761] & ~in[193]; 
    assign layer_0[6375] = ~(in[776] ^ in[673]); 
    assign layer_0[6376] = ~in[856]; 
    assign layer_0[6377] = in[485] ^ in[795]; 
    assign layer_0[6378] = 1'b0; 
    assign layer_0[6379] = ~(in[921] ^ in[974]); 
    assign layer_0[6380] = ~in[425] | (in[425] & in[461]); 
    assign layer_0[6381] = ~in[388] | (in[356] & in[388]); 
    assign layer_0[6382] = ~(in[452] ^ in[753]); 
    assign layer_0[6383] = in[55]; 
    assign layer_0[6384] = in[747]; 
    assign layer_0[6385] = in[937] | in[936]; 
    assign layer_0[6386] = ~in[806]; 
    assign layer_0[6387] = in[597] ^ in[262]; 
    assign layer_0[6388] = in[632] & ~in[347]; 
    assign layer_0[6389] = in[646] & in[621]; 
    assign layer_0[6390] = ~in[852]; 
    assign layer_0[6391] = in[933]; 
    assign layer_0[6392] = in[250] ^ in[1016]; 
    assign layer_0[6393] = ~in[309] | (in[913] & in[309]); 
    assign layer_0[6394] = ~in[49]; 
    assign layer_0[6395] = in[198]; 
    assign layer_0[6396] = ~(in[738] ^ in[675]); 
    assign layer_0[6397] = ~in[108] | (in[108] & in[529]); 
    assign layer_0[6398] = in[579] ^ in[949]; 
    assign layer_0[6399] = in[29] ^ in[506]; 
    assign layer_0[6400] = in[35] ^ in[277]; 
    assign layer_0[6401] = in[332] ^ in[837]; 
    assign layer_0[6402] = ~(in[717] & in[375]); 
    assign layer_0[6403] = ~in[160]; 
    assign layer_0[6404] = ~(in[796] ^ in[857]); 
    assign layer_0[6405] = in[105] & in[600]; 
    assign layer_0[6406] = in[749] ^ in[301]; 
    assign layer_0[6407] = in[1020] & ~in[1005]; 
    assign layer_0[6408] = ~in[690]; 
    assign layer_0[6409] = in[328] & in[604]; 
    assign layer_0[6410] = 1'b0; 
    assign layer_0[6411] = ~(in[824] & in[617]); 
    assign layer_0[6412] = in[207] ^ in[706]; 
    assign layer_0[6413] = in[918] ^ in[1001]; 
    assign layer_0[6414] = 1'b1; 
    assign layer_0[6415] = ~(in[496] | in[834]); 
    assign layer_0[6416] = in[420] ^ in[413]; 
    assign layer_0[6417] = in[963] | in[884]; 
    assign layer_0[6418] = ~(in[1019] | in[979]); 
    assign layer_0[6419] = ~(in[96] ^ in[958]); 
    assign layer_0[6420] = in[938] & ~in[590]; 
    assign layer_0[6421] = ~in[596]; 
    assign layer_0[6422] = ~(in[805] ^ in[173]); 
    assign layer_0[6423] = ~(in[874] | in[368]); 
    assign layer_0[6424] = ~(in[162] ^ in[349]); 
    assign layer_0[6425] = in[232] & in[465]; 
    assign layer_0[6426] = in[625] | in[943]; 
    assign layer_0[6427] = ~in[404] | (in[663] & in[404]); 
    assign layer_0[6428] = in[636] ^ in[756]; 
    assign layer_0[6429] = ~(in[472] ^ in[188]); 
    assign layer_0[6430] = ~(in[353] ^ in[898]); 
    assign layer_0[6431] = ~(in[532] ^ in[580]); 
    assign layer_0[6432] = in[573] ^ in[571]; 
    assign layer_0[6433] = in[1014] ^ in[914]; 
    assign layer_0[6434] = 1'b1; 
    assign layer_0[6435] = ~in[729] | (in[729] & in[260]); 
    assign layer_0[6436] = in[784] & ~in[953]; 
    assign layer_0[6437] = in[549] & ~in[387]; 
    assign layer_0[6438] = ~(in[4] ^ in[839]); 
    assign layer_0[6439] = in[212] & ~in[142]; 
    assign layer_0[6440] = in[655]; 
    assign layer_0[6441] = ~in[508]; 
    assign layer_0[6442] = in[748] & ~in[989]; 
    assign layer_0[6443] = ~(in[384] & in[401]); 
    assign layer_0[6444] = ~(in[616] ^ in[3]); 
    assign layer_0[6445] = ~in[586] | (in[586] & in[651]); 
    assign layer_0[6446] = in[919] ^ in[920]; 
    assign layer_0[6447] = in[650] ^ in[430]; 
    assign layer_0[6448] = in[835] ^ in[582]; 
    assign layer_0[6449] = ~(in[13] ^ in[885]); 
    assign layer_0[6450] = ~(in[714] | in[64]); 
    assign layer_0[6451] = ~in[923] | (in[923] & in[130]); 
    assign layer_0[6452] = ~in[307] | (in[307] & in[496]); 
    assign layer_0[6453] = ~in[345] | (in[869] & in[345]); 
    assign layer_0[6454] = in[510] & in[251]; 
    assign layer_0[6455] = in[966] & in[619]; 
    assign layer_0[6456] = ~in[935] | (in[935] & in[511]); 
    assign layer_0[6457] = in[298] | in[388]; 
    assign layer_0[6458] = ~(in[787] | in[241]); 
    assign layer_0[6459] = in[805]; 
    assign layer_0[6460] = ~(in[288] ^ in[246]); 
    assign layer_0[6461] = in[907] ^ in[4]; 
    assign layer_0[6462] = ~in[498]; 
    assign layer_0[6463] = 1'b1; 
    assign layer_0[6464] = ~in[651] | (in[987] & in[651]); 
    assign layer_0[6465] = in[957] ^ in[997]; 
    assign layer_0[6466] = ~in[971] | (in[971] & in[968]); 
    assign layer_0[6467] = ~(in[414] ^ in[711]); 
    assign layer_0[6468] = ~in[216] | (in[216] & in[5]); 
    assign layer_0[6469] = ~(in[461] | in[950]); 
    assign layer_0[6470] = in[628] ^ in[121]; 
    assign layer_0[6471] = ~(in[891] & in[598]); 
    assign layer_0[6472] = ~in[601]; 
    assign layer_0[6473] = in[396] & ~in[954]; 
    assign layer_0[6474] = in[340]; 
    assign layer_0[6475] = in[378] ^ in[325]; 
    assign layer_0[6476] = ~in[50]; 
    assign layer_0[6477] = ~(in[871] ^ in[463]); 
    assign layer_0[6478] = in[890] & ~in[208]; 
    assign layer_0[6479] = ~(in[996] ^ in[900]); 
    assign layer_0[6480] = ~(in[827] ^ in[387]); 
    assign layer_0[6481] = ~in[893] | (in[885] & in[893]); 
    assign layer_0[6482] = ~(in[757] ^ in[356]); 
    assign layer_0[6483] = in[306]; 
    assign layer_0[6484] = ~(in[886] ^ in[264]); 
    assign layer_0[6485] = in[967]; 
    assign layer_0[6486] = ~(in[87] | in[484]); 
    assign layer_0[6487] = ~(in[381] ^ in[644]); 
    assign layer_0[6488] = ~(in[413] ^ in[66]); 
    assign layer_0[6489] = in[584] ^ in[883]; 
    assign layer_0[6490] = in[63] ^ in[835]; 
    assign layer_0[6491] = in[474] | in[921]; 
    assign layer_0[6492] = ~(in[673] & in[416]); 
    assign layer_0[6493] = in[445] & ~in[278]; 
    assign layer_0[6494] = in[71] | in[760]; 
    assign layer_0[6495] = in[447] ^ in[28]; 
    assign layer_0[6496] = ~(in[979] ^ in[437]); 
    assign layer_0[6497] = ~(in[727] ^ in[733]); 
    assign layer_0[6498] = in[587] & ~in[749]; 
    assign layer_0[6499] = in[588] | in[940]; 
    assign layer_0[6500] = ~(in[371] & in[244]); 
    assign layer_0[6501] = in[867] ^ in[2]; 
    assign layer_0[6502] = ~(in[252] ^ in[587]); 
    assign layer_0[6503] = in[666] | in[173]; 
    assign layer_0[6504] = ~(in[1013] & in[495]); 
    assign layer_0[6505] = in[615] & in[682]; 
    assign layer_0[6506] = in[944] | in[984]; 
    assign layer_0[6507] = 1'b0; 
    assign layer_0[6508] = in[370] & ~in[874]; 
    assign layer_0[6509] = in[531]; 
    assign layer_0[6510] = ~(in[679] & in[217]); 
    assign layer_0[6511] = ~in[1016] | (in[357] & in[1016]); 
    assign layer_0[6512] = in[15] & ~in[233]; 
    assign layer_0[6513] = in[338] | in[987]; 
    assign layer_0[6514] = in[468] ^ in[116]; 
    assign layer_0[6515] = in[628]; 
    assign layer_0[6516] = ~(in[968] ^ in[458]); 
    assign layer_0[6517] = ~in[855]; 
    assign layer_0[6518] = ~(in[582] & in[950]); 
    assign layer_0[6519] = in[77] & ~in[870]; 
    assign layer_0[6520] = in[744]; 
    assign layer_0[6521] = in[782] | in[829]; 
    assign layer_0[6522] = in[807] & ~in[969]; 
    assign layer_0[6523] = ~in[41]; 
    assign layer_0[6524] = in[362] & ~in[79]; 
    assign layer_0[6525] = in[581] ^ in[564]; 
    assign layer_0[6526] = in[252] & in[424]; 
    assign layer_0[6527] = ~in[939]; 
    assign layer_0[6528] = ~in[85]; 
    assign layer_0[6529] = ~in[534]; 
    assign layer_0[6530] = 1'b1; 
    assign layer_0[6531] = ~in[851] | (in[851] & in[1015]); 
    assign layer_0[6532] = in[387] & in[9]; 
    assign layer_0[6533] = ~(in[316] ^ in[641]); 
    assign layer_0[6534] = ~(in[492] | in[995]); 
    assign layer_0[6535] = ~(in[517] | in[590]); 
    assign layer_0[6536] = in[885] ^ in[936]; 
    assign layer_0[6537] = in[724] & in[12]; 
    assign layer_0[6538] = ~(in[446] ^ in[443]); 
    assign layer_0[6539] = in[6] & in[660]; 
    assign layer_0[6540] = in[489] & in[554]; 
    assign layer_0[6541] = in[168] ^ in[852]; 
    assign layer_0[6542] = in[716] ^ in[264]; 
    assign layer_0[6543] = ~in[758] | (in[758] & in[693]); 
    assign layer_0[6544] = in[860] ^ in[627]; 
    assign layer_0[6545] = in[355] ^ in[233]; 
    assign layer_0[6546] = ~(in[926] ^ in[124]); 
    assign layer_0[6547] = ~(in[968] ^ in[133]); 
    assign layer_0[6548] = in[869] ^ in[587]; 
    assign layer_0[6549] = ~in[547] | (in[547] & in[530]); 
    assign layer_0[6550] = in[910] ^ in[60]; 
    assign layer_0[6551] = ~(in[699] ^ in[1001]); 
    assign layer_0[6552] = in[689] & ~in[730]; 
    assign layer_0[6553] = ~in[634]; 
    assign layer_0[6554] = in[12] ^ in[953]; 
    assign layer_0[6555] = in[294] ^ in[621]; 
    assign layer_0[6556] = ~in[653]; 
    assign layer_0[6557] = in[537]; 
    assign layer_0[6558] = in[900] & ~in[567]; 
    assign layer_0[6559] = ~(in[748] ^ in[637]); 
    assign layer_0[6560] = ~in[550] | (in[550] & in[301]); 
    assign layer_0[6561] = in[833] ^ in[703]; 
    assign layer_0[6562] = ~in[401] | (in[401] & in[772]); 
    assign layer_0[6563] = in[690] & ~in[499]; 
    assign layer_0[6564] = ~(in[793] ^ in[247]); 
    assign layer_0[6565] = ~(in[905] ^ in[601]); 
    assign layer_0[6566] = ~(in[460] ^ in[156]); 
    assign layer_0[6567] = in[648] & ~in[853]; 
    assign layer_0[6568] = in[804] ^ in[251]; 
    assign layer_0[6569] = ~(in[839] ^ in[837]); 
    assign layer_0[6570] = ~in[275]; 
    assign layer_0[6571] = ~(in[450] | in[129]); 
    assign layer_0[6572] = ~in[227] | (in[227] & in[916]); 
    assign layer_0[6573] = in[921] ^ in[339]; 
    assign layer_0[6574] = ~(in[705] ^ in[47]); 
    assign layer_0[6575] = ~(in[385] ^ in[834]); 
    assign layer_0[6576] = ~(in[536] & in[538]); 
    assign layer_0[6577] = in[646] & ~in[660]; 
    assign layer_0[6578] = in[291] | in[194]; 
    assign layer_0[6579] = in[857] | in[237]; 
    assign layer_0[6580] = in[623]; 
    assign layer_0[6581] = in[843] ^ in[704]; 
    assign layer_0[6582] = in[682] | in[447]; 
    assign layer_0[6583] = ~in[484]; 
    assign layer_0[6584] = ~(in[533] ^ in[522]); 
    assign layer_0[6585] = in[577] | in[129]; 
    assign layer_0[6586] = ~in[277] | (in[277] & in[843]); 
    assign layer_0[6587] = ~(in[210] ^ in[86]); 
    assign layer_0[6588] = ~in[454]; 
    assign layer_0[6589] = in[700]; 
    assign layer_0[6590] = ~(in[535] ^ in[588]); 
    assign layer_0[6591] = in[533] & ~in[987]; 
    assign layer_0[6592] = in[555]; 
    assign layer_0[6593] = ~in[389] | (in[999] & in[389]); 
    assign layer_0[6594] = ~(in[284] & in[311]); 
    assign layer_0[6595] = in[570] ^ in[950]; 
    assign layer_0[6596] = in[354] & ~in[742]; 
    assign layer_0[6597] = in[132] ^ in[724]; 
    assign layer_0[6598] = ~(in[676] ^ in[552]); 
    assign layer_0[6599] = in[873] ^ in[964]; 
    assign layer_0[6600] = in[8] & in[477]; 
    assign layer_0[6601] = in[330] & ~in[1019]; 
    assign layer_0[6602] = ~(in[275] ^ in[701]); 
    assign layer_0[6603] = ~(in[733] & in[333]); 
    assign layer_0[6604] = in[77] ^ in[803]; 
    assign layer_0[6605] = ~in[877]; 
    assign layer_0[6606] = ~(in[969] & in[936]); 
    assign layer_0[6607] = ~(in[593] | in[619]); 
    assign layer_0[6608] = in[649]; 
    assign layer_0[6609] = ~(in[920] ^ in[905]); 
    assign layer_0[6610] = ~(in[627] ^ in[641]); 
    assign layer_0[6611] = ~(in[61] ^ in[691]); 
    assign layer_0[6612] = in[852]; 
    assign layer_0[6613] = in[891] ^ in[551]; 
    assign layer_0[6614] = ~in[453] | (in[870] & in[453]); 
    assign layer_0[6615] = ~(in[348] & in[539]); 
    assign layer_0[6616] = ~(in[572] ^ in[448]); 
    assign layer_0[6617] = ~in[170] | (in[301] & in[170]); 
    assign layer_0[6618] = ~(in[294] | in[407]); 
    assign layer_0[6619] = in[985] ^ in[261]; 
    assign layer_0[6620] = in[701]; 
    assign layer_0[6621] = in[469] ^ in[108]; 
    assign layer_0[6622] = ~in[117]; 
    assign layer_0[6623] = ~in[748] | (in[748] & in[765]); 
    assign layer_0[6624] = in[923] | in[822]; 
    assign layer_0[6625] = in[49] ^ in[867]; 
    assign layer_0[6626] = ~(in[440] ^ in[333]); 
    assign layer_0[6627] = in[402] ^ in[915]; 
    assign layer_0[6628] = in[536] ^ in[725]; 
    assign layer_0[6629] = in[731] ^ in[692]; 
    assign layer_0[6630] = in[936] ^ in[276]; 
    assign layer_0[6631] = ~(in[885] ^ in[698]); 
    assign layer_0[6632] = in[918]; 
    assign layer_0[6633] = ~in[654]; 
    assign layer_0[6634] = in[565] & in[836]; 
    assign layer_0[6635] = in[936] ^ in[937]; 
    assign layer_0[6636] = ~(in[492] | in[719]); 
    assign layer_0[6637] = in[264] ^ in[322]; 
    assign layer_0[6638] = in[157] | in[555]; 
    assign layer_0[6639] = in[284] | in[611]; 
    assign layer_0[6640] = ~(in[775] ^ in[244]); 
    assign layer_0[6641] = in[741] & ~in[759]; 
    assign layer_0[6642] = in[744] ^ in[585]; 
    assign layer_0[6643] = 1'b1; 
    assign layer_0[6644] = in[518] ^ in[968]; 
    assign layer_0[6645] = ~in[267]; 
    assign layer_0[6646] = ~in[631] | (in[631] & in[732]); 
    assign layer_0[6647] = ~in[51] | (in[796] & in[51]); 
    assign layer_0[6648] = in[666] | in[858]; 
    assign layer_0[6649] = in[423] & ~in[513]; 
    assign layer_0[6650] = ~(in[435] ^ in[322]); 
    assign layer_0[6651] = ~(in[4] | in[1016]); 
    assign layer_0[6652] = ~(in[822] ^ in[195]); 
    assign layer_0[6653] = in[954]; 
    assign layer_0[6654] = in[694] & ~in[96]; 
    assign layer_0[6655] = in[1013]; 
    assign layer_0[6656] = ~(in[520] | in[875]); 
    assign layer_0[6657] = ~in[818] | (in[818] & in[221]); 
    assign layer_0[6658] = ~(in[709] ^ in[628]); 
    assign layer_0[6659] = 1'b0; 
    assign layer_0[6660] = ~(in[125] ^ in[1001]); 
    assign layer_0[6661] = in[638]; 
    assign layer_0[6662] = ~(in[386] ^ in[904]); 
    assign layer_0[6663] = ~(in[871] ^ in[859]); 
    assign layer_0[6664] = ~(in[35] ^ in[242]); 
    assign layer_0[6665] = ~(in[868] | in[872]); 
    assign layer_0[6666] = in[760] | in[572]; 
    assign layer_0[6667] = ~in[346]; 
    assign layer_0[6668] = in[868]; 
    assign layer_0[6669] = ~in[802] | (in[1011] & in[802]); 
    assign layer_0[6670] = ~(in[433] | in[471]); 
    assign layer_0[6671] = in[760] & ~in[891]; 
    assign layer_0[6672] = in[80] ^ in[138]; 
    assign layer_0[6673] = ~in[488] | (in[408] & in[488]); 
    assign layer_0[6674] = in[798]; 
    assign layer_0[6675] = ~in[348]; 
    assign layer_0[6676] = ~(in[754] | in[928]); 
    assign layer_0[6677] = ~in[917] | (in[917] & in[883]); 
    assign layer_0[6678] = ~in[724] | (in[724] & in[763]); 
    assign layer_0[6679] = ~(in[232] | in[322]); 
    assign layer_0[6680] = in[920] & in[41]; 
    assign layer_0[6681] = ~(in[498] ^ in[127]); 
    assign layer_0[6682] = ~(in[126] ^ in[190]); 
    assign layer_0[6683] = ~in[94]; 
    assign layer_0[6684] = in[211] & in[267]; 
    assign layer_0[6685] = ~(in[973] ^ in[896]); 
    assign layer_0[6686] = in[563]; 
    assign layer_0[6687] = in[1012] & ~in[664]; 
    assign layer_0[6688] = in[718]; 
    assign layer_0[6689] = ~(in[117] & in[195]); 
    assign layer_0[6690] = ~in[357] | (in[61] & in[357]); 
    assign layer_0[6691] = ~(in[413] ^ in[857]); 
    assign layer_0[6692] = in[857] ^ in[1021]; 
    assign layer_0[6693] = ~in[968] | (in[968] & in[994]); 
    assign layer_0[6694] = ~in[467] | (in[707] & in[467]); 
    assign layer_0[6695] = ~in[81]; 
    assign layer_0[6696] = ~in[670]; 
    assign layer_0[6697] = in[610] | in[398]; 
    assign layer_0[6698] = in[77] ^ in[295]; 
    assign layer_0[6699] = in[538] ^ in[900]; 
    assign layer_0[6700] = ~(in[184] & in[480]); 
    assign layer_0[6701] = ~(in[264] & in[62]); 
    assign layer_0[6702] = ~(in[429] ^ in[565]); 
    assign layer_0[6703] = in[520] ^ in[522]; 
    assign layer_0[6704] = ~in[857]; 
    assign layer_0[6705] = in[483] ^ in[905]; 
    assign layer_0[6706] = ~in[237] | (in[237] & in[1023]); 
    assign layer_0[6707] = in[615] ^ in[333]; 
    assign layer_0[6708] = in[417] & ~in[474]; 
    assign layer_0[6709] = in[186] & in[837]; 
    assign layer_0[6710] = ~in[947]; 
    assign layer_0[6711] = ~(in[346] & in[166]); 
    assign layer_0[6712] = ~(in[536] & in[28]); 
    assign layer_0[6713] = ~in[379] | (in[379] & in[848]); 
    assign layer_0[6714] = ~(in[571] | in[297]); 
    assign layer_0[6715] = in[949] ^ in[919]; 
    assign layer_0[6716] = in[1020] | in[449]; 
    assign layer_0[6717] = in[564]; 
    assign layer_0[6718] = in[99] ^ in[952]; 
    assign layer_0[6719] = in[872] ^ in[991]; 
    assign layer_0[6720] = ~(in[638] ^ in[748]); 
    assign layer_0[6721] = in[852]; 
    assign layer_0[6722] = in[595] & ~in[581]; 
    assign layer_0[6723] = in[220] ^ in[931]; 
    assign layer_0[6724] = in[956] & ~in[826]; 
    assign layer_0[6725] = ~(in[886] ^ in[616]); 
    assign layer_0[6726] = ~in[635]; 
    assign layer_0[6727] = ~in[507] | (in[811] & in[507]); 
    assign layer_0[6728] = ~in[21] | (in[256] & in[21]); 
    assign layer_0[6729] = ~in[469] | (in[469] & in[939]); 
    assign layer_0[6730] = in[211]; 
    assign layer_0[6731] = ~(in[842] ^ in[934]); 
    assign layer_0[6732] = in[902] & ~in[807]; 
    assign layer_0[6733] = ~(in[621] | in[593]); 
    assign layer_0[6734] = in[82] ^ in[45]; 
    assign layer_0[6735] = in[623] & ~in[733]; 
    assign layer_0[6736] = in[39] | in[961]; 
    assign layer_0[6737] = ~(in[769] | in[8]); 
    assign layer_0[6738] = in[684]; 
    assign layer_0[6739] = ~in[276] | (in[276] & in[852]); 
    assign layer_0[6740] = in[150] ^ in[73]; 
    assign layer_0[6741] = ~(in[73] ^ in[334]); 
    assign layer_0[6742] = in[897] ^ in[703]; 
    assign layer_0[6743] = in[666]; 
    assign layer_0[6744] = ~(in[129] & in[164]); 
    assign layer_0[6745] = in[759] & ~in[918]; 
    assign layer_0[6746] = in[773] ^ in[204]; 
    assign layer_0[6747] = in[414] & ~in[733]; 
    assign layer_0[6748] = ~(in[233] ^ in[777]); 
    assign layer_0[6749] = in[33] & ~in[803]; 
    assign layer_0[6750] = ~(in[141] ^ in[301]); 
    assign layer_0[6751] = in[806]; 
    assign layer_0[6752] = in[445] ^ in[280]; 
    assign layer_0[6753] = ~(in[1016] ^ in[260]); 
    assign layer_0[6754] = ~in[280] | (in[280] & in[550]); 
    assign layer_0[6755] = in[205] ^ in[625]; 
    assign layer_0[6756] = ~(in[605] & in[215]); 
    assign layer_0[6757] = ~(in[516] ^ in[306]); 
    assign layer_0[6758] = ~(in[276] ^ in[113]); 
    assign layer_0[6759] = 1'b0; 
    assign layer_0[6760] = in[476] ^ in[731]; 
    assign layer_0[6761] = in[971] & ~in[268]; 
    assign layer_0[6762] = ~in[471] | (in[471] & in[741]); 
    assign layer_0[6763] = ~in[933] | (in[933] & in[457]); 
    assign layer_0[6764] = ~in[160] | (in[160] & in[1019]); 
    assign layer_0[6765] = 1'b1; 
    assign layer_0[6766] = ~(in[486] ^ in[552]); 
    assign layer_0[6767] = ~in[51] | (in[51] & in[33]); 
    assign layer_0[6768] = in[82]; 
    assign layer_0[6769] = ~(in[389] | in[895]); 
    assign layer_0[6770] = in[426]; 
    assign layer_0[6771] = in[689]; 
    assign layer_0[6772] = ~in[221]; 
    assign layer_0[6773] = ~(in[908] ^ in[98]); 
    assign layer_0[6774] = in[984] ^ in[985]; 
    assign layer_0[6775] = ~(in[854] ^ in[932]); 
    assign layer_0[6776] = ~in[440]; 
    assign layer_0[6777] = in[364] ^ in[964]; 
    assign layer_0[6778] = ~in[994] | (in[639] & in[994]); 
    assign layer_0[6779] = in[810] | in[35]; 
    assign layer_0[6780] = ~(in[364] ^ in[492]); 
    assign layer_0[6781] = in[1014]; 
    assign layer_0[6782] = ~in[974] | (in[974] & in[406]); 
    assign layer_0[6783] = ~(in[640] ^ in[619]); 
    assign layer_0[6784] = ~(in[694] ^ in[535]); 
    assign layer_0[6785] = ~(in[897] | in[990]); 
    assign layer_0[6786] = ~(in[312] & in[253]); 
    assign layer_0[6787] = ~(in[779] ^ in[493]); 
    assign layer_0[6788] = in[318]; 
    assign layer_0[6789] = in[319] ^ in[615]; 
    assign layer_0[6790] = in[868] ^ in[878]; 
    assign layer_0[6791] = ~in[881]; 
    assign layer_0[6792] = ~(in[867] & in[604]); 
    assign layer_0[6793] = in[509] & ~in[360]; 
    assign layer_0[6794] = in[29] & ~in[392]; 
    assign layer_0[6795] = in[871] | in[606]; 
    assign layer_0[6796] = ~(in[382] & in[428]); 
    assign layer_0[6797] = ~(in[172] ^ in[572]); 
    assign layer_0[6798] = in[390] & ~in[234]; 
    assign layer_0[6799] = in[507] & in[584]; 
    assign layer_0[6800] = ~in[302]; 
    assign layer_0[6801] = ~(in[283] & in[744]); 
    assign layer_0[6802] = in[631] & ~in[624]; 
    assign layer_0[6803] = ~in[19] | (in[995] & in[19]); 
    assign layer_0[6804] = in[885] & ~in[870]; 
    assign layer_0[6805] = in[215] & ~in[568]; 
    assign layer_0[6806] = ~in[676] | (in[676] & in[708]); 
    assign layer_0[6807] = in[945] | in[507]; 
    assign layer_0[6808] = ~in[889] | (in[950] & in[889]); 
    assign layer_0[6809] = in[1018] ^ in[522]; 
    assign layer_0[6810] = in[451] ^ in[338]; 
    assign layer_0[6811] = in[950] ^ in[793]; 
    assign layer_0[6812] = ~(in[589] ^ in[79]); 
    assign layer_0[6813] = ~in[8]; 
    assign layer_0[6814] = ~(in[284] & in[613]); 
    assign layer_0[6815] = ~(in[617] & in[404]); 
    assign layer_0[6816] = 1'b1; 
    assign layer_0[6817] = in[791] & ~in[255]; 
    assign layer_0[6818] = ~in[328] | (in[845] & in[328]); 
    assign layer_0[6819] = in[673] & in[600]; 
    assign layer_0[6820] = ~in[755]; 
    assign layer_0[6821] = ~in[938] | (in[938] & in[888]); 
    assign layer_0[6822] = ~(in[989] ^ in[972]); 
    assign layer_0[6823] = ~(in[744] & in[748]); 
    assign layer_0[6824] = ~(in[917] ^ in[611]); 
    assign layer_0[6825] = in[970] ^ in[807]; 
    assign layer_0[6826] = ~(in[318] ^ in[906]); 
    assign layer_0[6827] = in[447] ^ in[719]; 
    assign layer_0[6828] = in[30] & ~in[530]; 
    assign layer_0[6829] = in[35]; 
    assign layer_0[6830] = in[627] & ~in[690]; 
    assign layer_0[6831] = 1'b0; 
    assign layer_0[6832] = in[177] ^ in[322]; 
    assign layer_0[6833] = in[970] | in[716]; 
    assign layer_0[6834] = ~in[243]; 
    assign layer_0[6835] = ~in[245]; 
    assign layer_0[6836] = in[201] ^ in[924]; 
    assign layer_0[6837] = in[808] ^ in[396]; 
    assign layer_0[6838] = in[604] | in[1018]; 
    assign layer_0[6839] = ~(in[172] | in[179]); 
    assign layer_0[6840] = in[30] ^ in[20]; 
    assign layer_0[6841] = ~(in[722] | in[416]); 
    assign layer_0[6842] = in[505] & ~in[723]; 
    assign layer_0[6843] = in[555] & ~in[563]; 
    assign layer_0[6844] = in[228]; 
    assign layer_0[6845] = ~in[259] | (in[259] & in[458]); 
    assign layer_0[6846] = ~(in[597] & in[237]); 
    assign layer_0[6847] = ~in[407] | (in[629] & in[407]); 
    assign layer_0[6848] = ~(in[587] & in[998]); 
    assign layer_0[6849] = ~in[728]; 
    assign layer_0[6850] = ~(in[549] ^ in[520]); 
    assign layer_0[6851] = ~(in[13] ^ in[1017]); 
    assign layer_0[6852] = ~(in[277] | in[416]); 
    assign layer_0[6853] = in[620] & ~in[431]; 
    assign layer_0[6854] = ~(in[465] & in[445]); 
    assign layer_0[6855] = ~in[186] | (in[186] & in[37]); 
    assign layer_0[6856] = in[264] & ~in[45]; 
    assign layer_0[6857] = in[463] & ~in[236]; 
    assign layer_0[6858] = in[663] ^ in[20]; 
    assign layer_0[6859] = in[250]; 
    assign layer_0[6860] = ~(in[107] & in[394]); 
    assign layer_0[6861] = ~(in[745] ^ in[744]); 
    assign layer_0[6862] = ~(in[1017] ^ in[318]); 
    assign layer_0[6863] = in[227] & in[99]; 
    assign layer_0[6864] = in[928] ^ in[956]; 
    assign layer_0[6865] = ~(in[712] ^ in[402]); 
    assign layer_0[6866] = in[145] & in[719]; 
    assign layer_0[6867] = ~(in[504] & in[372]); 
    assign layer_0[6868] = in[978]; 
    assign layer_0[6869] = in[587] & ~in[916]; 
    assign layer_0[6870] = ~(in[553] ^ in[844]); 
    assign layer_0[6871] = in[886] ^ in[568]; 
    assign layer_0[6872] = ~in[152] | (in[152] & in[724]); 
    assign layer_0[6873] = ~(in[842] ^ in[337]); 
    assign layer_0[6874] = ~in[314] | (in[314] & in[387]); 
    assign layer_0[6875] = in[66] & in[489]; 
    assign layer_0[6876] = in[503]; 
    assign layer_0[6877] = ~in[632] | (in[632] & in[272]); 
    assign layer_0[6878] = ~(in[747] ^ in[275]); 
    assign layer_0[6879] = in[548] ^ in[563]; 
    assign layer_0[6880] = ~(in[253] | in[349]); 
    assign layer_0[6881] = in[253] & ~in[971]; 
    assign layer_0[6882] = in[1015] | in[937]; 
    assign layer_0[6883] = ~(in[856] ^ in[906]); 
    assign layer_0[6884] = ~in[596]; 
    assign layer_0[6885] = ~(in[542] | in[522]); 
    assign layer_0[6886] = in[628] ^ in[683]; 
    assign layer_0[6887] = ~(in[62] ^ in[973]); 
    assign layer_0[6888] = in[952] ^ in[1001]; 
    assign layer_0[6889] = in[252] ^ in[202]; 
    assign layer_0[6890] = ~(in[380] ^ in[792]); 
    assign layer_0[6891] = ~(in[77] | in[563]); 
    assign layer_0[6892] = ~in[217]; 
    assign layer_0[6893] = in[49] ^ in[637]; 
    assign layer_0[6894] = in[646] & ~in[259]; 
    assign layer_0[6895] = ~(in[949] | in[513]); 
    assign layer_0[6896] = in[94]; 
    assign layer_0[6897] = in[611]; 
    assign layer_0[6898] = ~in[585]; 
    assign layer_0[6899] = ~in[9] | (in[9] & in[929]); 
    assign layer_0[6900] = in[986] & ~in[335]; 
    assign layer_0[6901] = in[120] ^ in[656]; 
    assign layer_0[6902] = ~in[537]; 
    assign layer_0[6903] = in[423] & in[95]; 
    assign layer_0[6904] = in[478]; 
    assign layer_0[6905] = ~in[64]; 
    assign layer_0[6906] = in[926] ^ in[811]; 
    assign layer_0[6907] = in[789] | in[697]; 
    assign layer_0[6908] = in[385] & ~in[855]; 
    assign layer_0[6909] = ~(in[911] ^ in[75]); 
    assign layer_0[6910] = in[859] ^ in[614]; 
    assign layer_0[6911] = in[28] & in[521]; 
    assign layer_0[6912] = in[284] | in[871]; 
    assign layer_0[6913] = ~(in[740] ^ in[682]); 
    assign layer_0[6914] = in[201] | in[718]; 
    assign layer_0[6915] = ~in[231] | (in[231] & in[435]); 
    assign layer_0[6916] = 1'b0; 
    assign layer_0[6917] = in[107] | in[899]; 
    assign layer_0[6918] = ~(in[12] & in[348]); 
    assign layer_0[6919] = ~(in[795] ^ in[882]); 
    assign layer_0[6920] = in[567] & ~in[61]; 
    assign layer_0[6921] = in[509] ^ in[649]; 
    assign layer_0[6922] = in[292] ^ in[392]; 
    assign layer_0[6923] = ~in[9]; 
    assign layer_0[6924] = ~in[997] | (in[909] & in[997]); 
    assign layer_0[6925] = ~in[852] | (in[852] & in[266]); 
    assign layer_0[6926] = in[886] | in[822]; 
    assign layer_0[6927] = ~in[251]; 
    assign layer_0[6928] = ~in[903]; 
    assign layer_0[6929] = in[413]; 
    assign layer_0[6930] = in[1001]; 
    assign layer_0[6931] = in[579]; 
    assign layer_0[6932] = in[747] & ~in[990]; 
    assign layer_0[6933] = in[863] | in[846]; 
    assign layer_0[6934] = ~in[910] | (in[790] & in[910]); 
    assign layer_0[6935] = ~(in[145] | in[827]); 
    assign layer_0[6936] = in[195] & in[293]; 
    assign layer_0[6937] = ~in[666] | (in[666] & in[981]); 
    assign layer_0[6938] = ~in[75] | (in[692] & in[75]); 
    assign layer_0[6939] = in[7] & ~in[869]; 
    assign layer_0[6940] = ~in[608]; 
    assign layer_0[6941] = in[968] ^ in[483]; 
    assign layer_0[6942] = ~(in[312] ^ in[87]); 
    assign layer_0[6943] = ~in[891] | (in[508] & in[891]); 
    assign layer_0[6944] = in[883] | in[869]; 
    assign layer_0[6945] = in[688] ^ in[652]; 
    assign layer_0[6946] = ~in[630]; 
    assign layer_0[6947] = in[953] ^ in[130]; 
    assign layer_0[6948] = in[790]; 
    assign layer_0[6949] = in[679] ^ in[612]; 
    assign layer_0[6950] = ~(in[82] & in[381]); 
    assign layer_0[6951] = in[253]; 
    assign layer_0[6952] = in[851]; 
    assign layer_0[6953] = ~(in[686] ^ in[548]); 
    assign layer_0[6954] = ~(in[317] ^ in[599]); 
    assign layer_0[6955] = ~(in[852] ^ in[988]); 
    assign layer_0[6956] = in[277] | in[580]; 
    assign layer_0[6957] = 1'b0; 
    assign layer_0[6958] = in[549] & ~in[473]; 
    assign layer_0[6959] = ~(in[612] ^ in[446]); 
    assign layer_0[6960] = ~in[298] | (in[499] & in[298]); 
    assign layer_0[6961] = ~(in[262] ^ in[718]); 
    assign layer_0[6962] = in[955] ^ in[971]; 
    assign layer_0[6963] = in[892] | in[856]; 
    assign layer_0[6964] = ~in[570] | (in[917] & in[570]); 
    assign layer_0[6965] = in[231] & in[597]; 
    assign layer_0[6966] = in[762] ^ in[885]; 
    assign layer_0[6967] = in[617] & in[5]; 
    assign layer_0[6968] = in[61] ^ in[189]; 
    assign layer_0[6969] = ~in[556]; 
    assign layer_0[6970] = ~in[951] | (in[951] & in[862]); 
    assign layer_0[6971] = ~in[86] | (in[86] & in[539]); 
    assign layer_0[6972] = in[355]; 
    assign layer_0[6973] = in[96] ^ in[733]; 
    assign layer_0[6974] = ~(in[261] ^ in[786]); 
    assign layer_0[6975] = in[838] ^ in[28]; 
    assign layer_0[6976] = in[508] | in[224]; 
    assign layer_0[6977] = ~(in[433] | in[777]); 
    assign layer_0[6978] = in[934]; 
    assign layer_0[6979] = ~(in[841] ^ in[822]); 
    assign layer_0[6980] = ~(in[776] & in[297]); 
    assign layer_0[6981] = ~(in[556] ^ in[700]); 
    assign layer_0[6982] = in[325] & in[267]; 
    assign layer_0[6983] = ~(in[69] ^ in[704]); 
    assign layer_0[6984] = ~(in[814] | in[911]); 
    assign layer_0[6985] = in[920] & ~in[852]; 
    assign layer_0[6986] = in[692] & ~in[571]; 
    assign layer_0[6987] = in[664] ^ in[426]; 
    assign layer_0[6988] = in[413] ^ in[685]; 
    assign layer_0[6989] = ~(in[472] & in[99]); 
    assign layer_0[6990] = ~(in[630] & in[1013]); 
    assign layer_0[6991] = in[607] & ~in[241]; 
    assign layer_0[6992] = ~(in[605] & in[298]); 
    assign layer_0[6993] = ~(in[690] ^ in[126]); 
    assign layer_0[6994] = ~in[704]; 
    assign layer_0[6995] = ~(in[871] ^ in[724]); 
    assign layer_0[6996] = 1'b0; 
    assign layer_0[6997] = ~(in[671] ^ in[380]); 
    assign layer_0[6998] = ~(in[731] ^ in[701]); 
    assign layer_0[6999] = ~in[267]; 
    assign layer_0[7000] = in[457] | in[80]; 
    assign layer_0[7001] = ~(in[581] ^ in[533]); 
    assign layer_0[7002] = in[104] & in[177]; 
    assign layer_0[7003] = ~(in[325] | in[626]); 
    assign layer_0[7004] = ~in[431]; 
    assign layer_0[7005] = ~(in[869] | in[881]); 
    assign layer_0[7006] = in[524] & ~in[919]; 
    assign layer_0[7007] = ~in[263] | (in[263] & in[789]); 
    assign layer_0[7008] = ~(in[477] ^ in[967]); 
    assign layer_0[7009] = in[618] ^ in[762]; 
    assign layer_0[7010] = in[333]; 
    assign layer_0[7011] = ~in[655]; 
    assign layer_0[7012] = in[938] & ~in[898]; 
    assign layer_0[7013] = in[771]; 
    assign layer_0[7014] = in[765]; 
    assign layer_0[7015] = in[292] ^ in[905]; 
    assign layer_0[7016] = ~in[156] | (in[757] & in[156]); 
    assign layer_0[7017] = ~(in[935] ^ in[508]); 
    assign layer_0[7018] = in[920] ^ in[905]; 
    assign layer_0[7019] = ~(in[645] | in[623]); 
    assign layer_0[7020] = in[362] ^ in[808]; 
    assign layer_0[7021] = in[438] ^ in[951]; 
    assign layer_0[7022] = ~in[469]; 
    assign layer_0[7023] = in[300] | in[570]; 
    assign layer_0[7024] = ~in[665] | (in[665] & in[245]); 
    assign layer_0[7025] = ~(in[981] ^ in[955]); 
    assign layer_0[7026] = ~in[676] | (in[732] & in[676]); 
    assign layer_0[7027] = in[100]; 
    assign layer_0[7028] = in[566]; 
    assign layer_0[7029] = in[103] | in[108]; 
    assign layer_0[7030] = ~in[867]; 
    assign layer_0[7031] = ~(in[645] ^ in[56]); 
    assign layer_0[7032] = in[764]; 
    assign layer_0[7033] = in[888] ^ in[859]; 
    assign layer_0[7034] = in[440] & ~in[998]; 
    assign layer_0[7035] = ~(in[617] & in[450]); 
    assign layer_0[7036] = in[445] ^ in[581]; 
    assign layer_0[7037] = ~in[445]; 
    assign layer_0[7038] = in[180] & in[324]; 
    assign layer_0[7039] = in[531] ^ in[460]; 
    assign layer_0[7040] = ~(in[539] ^ in[740]); 
    assign layer_0[7041] = in[753]; 
    assign layer_0[7042] = ~(in[805] ^ in[824]); 
    assign layer_0[7043] = 1'b1; 
    assign layer_0[7044] = ~in[312]; 
    assign layer_0[7045] = ~(in[760] & in[203]); 
    assign layer_0[7046] = ~in[842] | (in[842] & in[519]); 
    assign layer_0[7047] = ~(in[315] & in[743]); 
    assign layer_0[7048] = in[483] ^ in[673]; 
    assign layer_0[7049] = ~in[481] | (in[589] & in[481]); 
    assign layer_0[7050] = in[970] | in[406]; 
    assign layer_0[7051] = ~(in[610] ^ in[621]); 
    assign layer_0[7052] = in[874]; 
    assign layer_0[7053] = ~in[334]; 
    assign layer_0[7054] = ~(in[61] | in[1016]); 
    assign layer_0[7055] = in[193] ^ in[732]; 
    assign layer_0[7056] = ~in[587]; 
    assign layer_0[7057] = ~(in[141] & in[728]); 
    assign layer_0[7058] = ~in[930]; 
    assign layer_0[7059] = ~(in[844] ^ in[626]); 
    assign layer_0[7060] = ~in[674] | (in[80] & in[674]); 
    assign layer_0[7061] = ~in[681]; 
    assign layer_0[7062] = ~in[679]; 
    assign layer_0[7063] = in[389] ^ in[864]; 
    assign layer_0[7064] = ~(in[955] ^ in[979]); 
    assign layer_0[7065] = ~(in[922] & in[627]); 
    assign layer_0[7066] = in[445]; 
    assign layer_0[7067] = ~(in[673] ^ in[79]); 
    assign layer_0[7068] = ~in[21]; 
    assign layer_0[7069] = in[61] & in[596]; 
    assign layer_0[7070] = in[386] & ~in[692]; 
    assign layer_0[7071] = in[642]; 
    assign layer_0[7072] = in[473] & ~in[519]; 
    assign layer_0[7073] = ~in[387] | (in[387] & in[587]); 
    assign layer_0[7074] = in[12] & ~in[541]; 
    assign layer_0[7075] = in[667]; 
    assign layer_0[7076] = ~in[336] | (in[141] & in[336]); 
    assign layer_0[7077] = in[188] ^ in[961]; 
    assign layer_0[7078] = ~(in[667] ^ in[808]); 
    assign layer_0[7079] = ~(in[79] ^ in[52]); 
    assign layer_0[7080] = ~in[898]; 
    assign layer_0[7081] = in[123] ^ in[597]; 
    assign layer_0[7082] = in[477] | in[965]; 
    assign layer_0[7083] = ~in[399] | (in[399] & in[967]); 
    assign layer_0[7084] = in[473]; 
    assign layer_0[7085] = ~in[268] | (in[48] & in[268]); 
    assign layer_0[7086] = in[806] ^ in[964]; 
    assign layer_0[7087] = in[568] ^ in[863]; 
    assign layer_0[7088] = ~in[218]; 
    assign layer_0[7089] = in[854] | in[259]; 
    assign layer_0[7090] = ~in[914]; 
    assign layer_0[7091] = ~(in[606] ^ in[629]); 
    assign layer_0[7092] = ~in[953]; 
    assign layer_0[7093] = ~(in[789] & in[695]); 
    assign layer_0[7094] = ~(in[873] ^ in[937]); 
    assign layer_0[7095] = in[485] ^ in[93]; 
    assign layer_0[7096] = in[642] & ~in[589]; 
    assign layer_0[7097] = ~(in[660] ^ in[571]); 
    assign layer_0[7098] = ~(in[624] | in[773]); 
    assign layer_0[7099] = ~(in[476] ^ in[876]); 
    assign layer_0[7100] = ~(in[988] & in[963]); 
    assign layer_0[7101] = in[807] ^ in[953]; 
    assign layer_0[7102] = ~in[372] | (in[372] & in[890]); 
    assign layer_0[7103] = in[871] & in[639]; 
    assign layer_0[7104] = in[921]; 
    assign layer_0[7105] = ~(in[394] | in[945]); 
    assign layer_0[7106] = in[526] ^ in[943]; 
    assign layer_0[7107] = ~in[424] | (in[424] & in[954]); 
    assign layer_0[7108] = in[265]; 
    assign layer_0[7109] = in[411] ^ in[688]; 
    assign layer_0[7110] = in[85] ^ in[940]; 
    assign layer_0[7111] = ~(in[124] & in[533]); 
    assign layer_0[7112] = in[177] ^ in[649]; 
    assign layer_0[7113] = ~(in[630] | in[517]); 
    assign layer_0[7114] = ~in[597]; 
    assign layer_0[7115] = in[220] ^ in[552]; 
    assign layer_0[7116] = ~in[165] | (in[691] & in[165]); 
    assign layer_0[7117] = ~in[574] | (in[911] & in[574]); 
    assign layer_0[7118] = in[405]; 
    assign layer_0[7119] = ~(in[952] ^ in[707]); 
    assign layer_0[7120] = ~in[659] | (in[659] & in[774]); 
    assign layer_0[7121] = in[300]; 
    assign layer_0[7122] = in[826]; 
    assign layer_0[7123] = in[209] & ~in[276]; 
    assign layer_0[7124] = in[637] | in[88]; 
    assign layer_0[7125] = in[262]; 
    assign layer_0[7126] = ~(in[579] ^ in[602]); 
    assign layer_0[7127] = ~(in[693] | in[480]); 
    assign layer_0[7128] = ~(in[595] ^ in[983]); 
    assign layer_0[7129] = in[692] ^ in[551]; 
    assign layer_0[7130] = in[193] & in[594]; 
    assign layer_0[7131] = ~in[969]; 
    assign layer_0[7132] = in[966]; 
    assign layer_0[7133] = in[933] & ~in[683]; 
    assign layer_0[7134] = ~(in[911] | in[94]); 
    assign layer_0[7135] = in[209]; 
    assign layer_0[7136] = ~in[707]; 
    assign layer_0[7137] = ~in[584] | (in[333] & in[584]); 
    assign layer_0[7138] = in[113]; 
    assign layer_0[7139] = ~(in[174] | in[0]); 
    assign layer_0[7140] = ~in[615] | (in[615] & in[731]); 
    assign layer_0[7141] = in[550] | in[844]; 
    assign layer_0[7142] = in[663]; 
    assign layer_0[7143] = ~(in[859] ^ in[519]); 
    assign layer_0[7144] = ~in[140]; 
    assign layer_0[7145] = in[889] | in[194]; 
    assign layer_0[7146] = ~(in[365] & in[296]); 
    assign layer_0[7147] = ~(in[673] | in[227]); 
    assign layer_0[7148] = ~(in[383] | in[994]); 
    assign layer_0[7149] = ~in[674]; 
    assign layer_0[7150] = ~(in[843] ^ in[778]); 
    assign layer_0[7151] = ~(in[932] ^ in[945]); 
    assign layer_0[7152] = in[212] ^ in[929]; 
    assign layer_0[7153] = ~(in[648] ^ in[679]); 
    assign layer_0[7154] = in[706] & in[901]; 
    assign layer_0[7155] = ~in[922]; 
    assign layer_0[7156] = in[867] & ~in[942]; 
    assign layer_0[7157] = ~in[907] | (in[900] & in[907]); 
    assign layer_0[7158] = ~(in[433] | in[4]); 
    assign layer_0[7159] = in[880]; 
    assign layer_0[7160] = in[349] ^ in[619]; 
    assign layer_0[7161] = ~(in[580] & in[74]); 
    assign layer_0[7162] = ~in[916] | (in[624] & in[916]); 
    assign layer_0[7163] = in[762]; 
    assign layer_0[7164] = in[802] & ~in[57]; 
    assign layer_0[7165] = in[714] & in[584]; 
    assign layer_0[7166] = ~(in[1019] | in[78]); 
    assign layer_0[7167] = in[266] | in[942]; 
    assign layer_0[7168] = ~in[376] | (in[998] & in[376]); 
    assign layer_0[7169] = ~(in[902] ^ in[970]); 
    assign layer_0[7170] = in[888] ^ in[856]; 
    assign layer_0[7171] = ~in[883] | (in[794] & in[883]); 
    assign layer_0[7172] = in[858] ^ in[820]; 
    assign layer_0[7173] = ~(in[675] ^ in[299]); 
    assign layer_0[7174] = ~(in[354] | in[997]); 
    assign layer_0[7175] = in[748]; 
    assign layer_0[7176] = in[538] & ~in[304]; 
    assign layer_0[7177] = ~(in[470] ^ in[3]); 
    assign layer_0[7178] = ~(in[950] | in[200]); 
    assign layer_0[7179] = ~in[303] | (in[303] & in[599]); 
    assign layer_0[7180] = ~in[931]; 
    assign layer_0[7181] = in[887] ^ in[668]; 
    assign layer_0[7182] = in[927] ^ in[310]; 
    assign layer_0[7183] = in[428] & in[902]; 
    assign layer_0[7184] = in[913] ^ in[931]; 
    assign layer_0[7185] = in[957] ^ in[1013]; 
    assign layer_0[7186] = ~(in[572] ^ in[417]); 
    assign layer_0[7187] = ~in[574]; 
    assign layer_0[7188] = 1'b0; 
    assign layer_0[7189] = 1'b1; 
    assign layer_0[7190] = ~in[646] | (in[564] & in[646]); 
    assign layer_0[7191] = in[568] & ~in[869]; 
    assign layer_0[7192] = ~in[967]; 
    assign layer_0[7193] = ~in[233]; 
    assign layer_0[7194] = ~(in[901] ^ in[810]); 
    assign layer_0[7195] = in[194] & ~in[951]; 
    assign layer_0[7196] = in[842] ^ in[620]; 
    assign layer_0[7197] = in[1013] | in[383]; 
    assign layer_0[7198] = in[109]; 
    assign layer_0[7199] = in[252] ^ in[364]; 
    assign layer_0[7200] = in[45] & in[546]; 
    assign layer_0[7201] = ~(in[920] ^ in[571]); 
    assign layer_0[7202] = in[727]; 
    assign layer_0[7203] = in[515] ^ in[252]; 
    assign layer_0[7204] = in[831] | in[1016]; 
    assign layer_0[7205] = ~(in[300] & in[508]); 
    assign layer_0[7206] = in[403] ^ in[1014]; 
    assign layer_0[7207] = in[935] & ~in[785]; 
    assign layer_0[7208] = in[469] & ~in[422]; 
    assign layer_0[7209] = in[466] ^ in[145]; 
    assign layer_0[7210] = ~in[582]; 
    assign layer_0[7211] = ~(in[935] ^ in[934]); 
    assign layer_0[7212] = ~in[323]; 
    assign layer_0[7213] = ~(in[600] ^ in[604]); 
    assign layer_0[7214] = in[366] ^ in[891]; 
    assign layer_0[7215] = in[376] & in[552]; 
    assign layer_0[7216] = in[35]; 
    assign layer_0[7217] = ~in[553] | (in[262] & in[553]); 
    assign layer_0[7218] = ~(in[519] ^ in[717]); 
    assign layer_0[7219] = ~(in[218] ^ in[223]); 
    assign layer_0[7220] = ~(in[916] ^ in[88]); 
    assign layer_0[7221] = ~(in[992] ^ in[13]); 
    assign layer_0[7222] = in[602] | in[969]; 
    assign layer_0[7223] = ~in[283]; 
    assign layer_0[7224] = in[855] & ~in[563]; 
    assign layer_0[7225] = in[122]; 
    assign layer_0[7226] = in[75] ^ in[862]; 
    assign layer_0[7227] = ~in[744] | (in[653] & in[744]); 
    assign layer_0[7228] = ~(in[935] & in[506]); 
    assign layer_0[7229] = ~(in[450] ^ in[833]); 
    assign layer_0[7230] = ~(in[263] ^ in[261]); 
    assign layer_0[7231] = ~(in[534] | in[322]); 
    assign layer_0[7232] = ~in[858]; 
    assign layer_0[7233] = ~(in[456] & in[8]); 
    assign layer_0[7234] = 1'b0; 
    assign layer_0[7235] = in[120] & in[82]; 
    assign layer_0[7236] = ~(in[966] ^ in[556]); 
    assign layer_0[7237] = ~in[512] | (in[764] & in[512]); 
    assign layer_0[7238] = in[846] | in[552]; 
    assign layer_0[7239] = ~in[297]; 
    assign layer_0[7240] = in[681] & in[8]; 
    assign layer_0[7241] = in[778]; 
    assign layer_0[7242] = ~(in[661] ^ in[873]); 
    assign layer_0[7243] = ~(in[999] | in[479]); 
    assign layer_0[7244] = 1'b0; 
    assign layer_0[7245] = in[62]; 
    assign layer_0[7246] = in[842] ^ in[884]; 
    assign layer_0[7247] = ~in[634]; 
    assign layer_0[7248] = in[906]; 
    assign layer_0[7249] = in[74] & ~in[734]; 
    assign layer_0[7250] = in[504]; 
    assign layer_0[7251] = ~(in[905] ^ in[920]); 
    assign layer_0[7252] = ~in[446]; 
    assign layer_0[7253] = ~in[389] | (in[389] & in[598]); 
    assign layer_0[7254] = ~(in[85] ^ in[562]); 
    assign layer_0[7255] = ~(in[808] ^ in[269]); 
    assign layer_0[7256] = ~in[888] | (in[888] & in[760]); 
    assign layer_0[7257] = in[889] ^ in[108]; 
    assign layer_0[7258] = in[63]; 
    assign layer_0[7259] = ~in[86] | (in[589] & in[86]); 
    assign layer_0[7260] = ~(in[417] & in[105]); 
    assign layer_0[7261] = in[302] & in[638]; 
    assign layer_0[7262] = in[2] | in[560]; 
    assign layer_0[7263] = in[210]; 
    assign layer_0[7264] = ~(in[891] ^ in[926]); 
    assign layer_0[7265] = ~in[604] | (in[477] & in[604]); 
    assign layer_0[7266] = in[1014] & ~in[477]; 
    assign layer_0[7267] = in[261]; 
    assign layer_0[7268] = ~(in[91] | in[785]); 
    assign layer_0[7269] = in[197]; 
    assign layer_0[7270] = in[481] & in[366]; 
    assign layer_0[7271] = ~(in[601] ^ in[859]); 
    assign layer_0[7272] = ~in[844]; 
    assign layer_0[7273] = in[18] | in[323]; 
    assign layer_0[7274] = in[364] ^ in[520]; 
    assign layer_0[7275] = ~(in[691] | in[161]); 
    assign layer_0[7276] = in[902] ^ in[888]; 
    assign layer_0[7277] = ~(in[986] | in[969]); 
    assign layer_0[7278] = ~in[556]; 
    assign layer_0[7279] = in[282] & ~in[827]; 
    assign layer_0[7280] = in[23]; 
    assign layer_0[7281] = in[713] ^ in[660]; 
    assign layer_0[7282] = in[708] & ~in[755]; 
    assign layer_0[7283] = in[739]; 
    assign layer_0[7284] = ~(in[392] & in[201]); 
    assign layer_0[7285] = ~in[265]; 
    assign layer_0[7286] = in[596] ^ in[724]; 
    assign layer_0[7287] = ~(in[623] ^ in[195]); 
    assign layer_0[7288] = ~in[446]; 
    assign layer_0[7289] = in[396] & ~in[515]; 
    assign layer_0[7290] = in[1001] ^ in[1000]; 
    assign layer_0[7291] = ~in[170] | (in[634] & in[170]); 
    assign layer_0[7292] = in[882]; 
    assign layer_0[7293] = ~(in[240] & in[283]); 
    assign layer_0[7294] = ~(in[59] ^ in[132]); 
    assign layer_0[7295] = ~(in[589] ^ in[938]); 
    assign layer_0[7296] = ~in[407]; 
    assign layer_0[7297] = in[367] ^ in[905]; 
    assign layer_0[7298] = ~(in[665] ^ in[582]); 
    assign layer_0[7299] = in[561]; 
    assign layer_0[7300] = ~(in[919] ^ in[102]); 
    assign layer_0[7301] = in[392] & ~in[899]; 
    assign layer_0[7302] = in[938] & in[892]; 
    assign layer_0[7303] = ~(in[97] ^ in[839]); 
    assign layer_0[7304] = ~in[551] | (in[540] & in[551]); 
    assign layer_0[7305] = ~(in[856] | in[783]); 
    assign layer_0[7306] = in[511] | in[615]; 
    assign layer_0[7307] = in[989] ^ in[547]; 
    assign layer_0[7308] = ~(in[676] & in[634]); 
    assign layer_0[7309] = ~in[713] | (in[713] & in[826]); 
    assign layer_0[7310] = in[423] & in[669]; 
    assign layer_0[7311] = ~(in[140] & in[851]); 
    assign layer_0[7312] = in[869] & ~in[924]; 
    assign layer_0[7313] = ~(in[349] ^ in[113]); 
    assign layer_0[7314] = ~in[62] | (in[572] & in[62]); 
    assign layer_0[7315] = ~in[673] | (in[673] & in[788]); 
    assign layer_0[7316] = ~(in[338] | in[764]); 
    assign layer_0[7317] = ~(in[793] | in[792]); 
    assign layer_0[7318] = in[741] ^ in[748]; 
    assign layer_0[7319] = in[921] ^ in[923]; 
    assign layer_0[7320] = ~in[773] | (in[65] & in[773]); 
    assign layer_0[7321] = ~in[129]; 
    assign layer_0[7322] = ~(in[146] | in[93]); 
    assign layer_0[7323] = ~(in[268] | in[703]); 
    assign layer_0[7324] = ~in[374]; 
    assign layer_0[7325] = in[281] & ~in[756]; 
    assign layer_0[7326] = in[984]; 
    assign layer_0[7327] = in[603] & ~in[477]; 
    assign layer_0[7328] = in[870] ^ in[851]; 
    assign layer_0[7329] = in[169] & in[56]; 
    assign layer_0[7330] = in[417] ^ in[855]; 
    assign layer_0[7331] = in[858] | in[78]; 
    assign layer_0[7332] = in[855] ^ in[824]; 
    assign layer_0[7333] = ~in[37] | (in[76] & in[37]); 
    assign layer_0[7334] = in[61] & ~in[786]; 
    assign layer_0[7335] = in[355] ^ in[211]; 
    assign layer_0[7336] = in[851] & ~in[933]; 
    assign layer_0[7337] = in[794] ^ in[676]; 
    assign layer_0[7338] = ~(in[877] ^ in[926]); 
    assign layer_0[7339] = in[602] ^ in[871]; 
    assign layer_0[7340] = ~in[805] | (in[805] & in[985]); 
    assign layer_0[7341] = in[226]; 
    assign layer_0[7342] = in[83]; 
    assign layer_0[7343] = in[761] ^ in[285]; 
    assign layer_0[7344] = in[438]; 
    assign layer_0[7345] = in[283] ^ in[808]; 
    assign layer_0[7346] = ~(in[980] ^ in[366]); 
    assign layer_0[7347] = ~in[252]; 
    assign layer_0[7348] = in[307] ^ in[969]; 
    assign layer_0[7349] = ~(in[972] ^ in[533]); 
    assign layer_0[7350] = in[11] & in[277]; 
    assign layer_0[7351] = in[417] & ~in[413]; 
    assign layer_0[7352] = in[502] | in[941]; 
    assign layer_0[7353] = ~(in[628] ^ in[616]); 
    assign layer_0[7354] = in[603] & ~in[526]; 
    assign layer_0[7355] = ~(in[630] & in[657]); 
    assign layer_0[7356] = ~(in[500] ^ in[948]); 
    assign layer_0[7357] = ~(in[980] & in[215]); 
    assign layer_0[7358] = in[970] ^ in[557]; 
    assign layer_0[7359] = in[365] & ~in[257]; 
    assign layer_0[7360] = in[68] | in[290]; 
    assign layer_0[7361] = in[770]; 
    assign layer_0[7362] = ~in[984]; 
    assign layer_0[7363] = in[668] ^ in[158]; 
    assign layer_0[7364] = in[139] ^ in[949]; 
    assign layer_0[7365] = ~in[699] | (in[355] & in[699]); 
    assign layer_0[7366] = 1'b1; 
    assign layer_0[7367] = ~(in[870] ^ in[902]); 
    assign layer_0[7368] = ~(in[129] ^ in[907]); 
    assign layer_0[7369] = ~(in[961] | in[450]); 
    assign layer_0[7370] = ~in[324]; 
    assign layer_0[7371] = ~in[263] | (in[263] & in[887]); 
    assign layer_0[7372] = in[74] ^ in[966]; 
    assign layer_0[7373] = ~(in[451] | in[882]); 
    assign layer_0[7374] = in[952] ^ in[897]; 
    assign layer_0[7375] = ~(in[522] ^ in[403]); 
    assign layer_0[7376] = in[225] & ~in[989]; 
    assign layer_0[7377] = in[895]; 
    assign layer_0[7378] = in[613] ^ in[265]; 
    assign layer_0[7379] = in[11]; 
    assign layer_0[7380] = in[887] ^ in[399]; 
    assign layer_0[7381] = in[838] ^ in[906]; 
    assign layer_0[7382] = in[903] ^ in[921]; 
    assign layer_0[7383] = ~(in[970] ^ in[969]); 
    assign layer_0[7384] = in[474] ^ in[763]; 
    assign layer_0[7385] = ~(in[950] & in[871]); 
    assign layer_0[7386] = in[666]; 
    assign layer_0[7387] = ~(in[437] | in[990]); 
    assign layer_0[7388] = ~(in[963] | in[1017]); 
    assign layer_0[7389] = in[689] | in[510]; 
    assign layer_0[7390] = ~(in[448] ^ in[1018]); 
    assign layer_0[7391] = in[850] & ~in[960]; 
    assign layer_0[7392] = in[580]; 
    assign layer_0[7393] = in[443] ^ in[586]; 
    assign layer_0[7394] = ~in[689] | (in[689] & in[461]); 
    assign layer_0[7395] = in[555] ^ in[284]; 
    assign layer_0[7396] = ~(in[386] ^ in[635]); 
    assign layer_0[7397] = ~(in[831] | in[553]); 
    assign layer_0[7398] = ~(in[29] ^ in[999]); 
    assign layer_0[7399] = ~(in[128] ^ in[445]); 
    assign layer_0[7400] = ~(in[591] ^ in[461]); 
    assign layer_0[7401] = in[221] & ~in[267]; 
    assign layer_0[7402] = ~(in[50] & in[461]); 
    assign layer_0[7403] = in[195] ^ in[220]; 
    assign layer_0[7404] = ~in[743] | (in[743] & in[1016]); 
    assign layer_0[7405] = in[697]; 
    assign layer_0[7406] = in[436] & in[854]; 
    assign layer_0[7407] = ~in[476] | (in[671] & in[476]); 
    assign layer_0[7408] = ~in[422]; 
    assign layer_0[7409] = ~(in[197] & in[719]); 
    assign layer_0[7410] = ~(in[968] ^ in[984]); 
    assign layer_0[7411] = ~in[644]; 
    assign layer_0[7412] = ~in[103] | (in[103] & in[420]); 
    assign layer_0[7413] = ~in[733]; 
    assign layer_0[7414] = in[685]; 
    assign layer_0[7415] = 1'b1; 
    assign layer_0[7416] = ~(in[191] & in[161]); 
    assign layer_0[7417] = ~(in[339] ^ in[587]); 
    assign layer_0[7418] = 1'b0; 
    assign layer_0[7419] = in[572] ^ in[499]; 
    assign layer_0[7420] = ~(in[596] ^ in[420]); 
    assign layer_0[7421] = ~(in[356] ^ in[793]); 
    assign layer_0[7422] = in[637] & in[635]; 
    assign layer_0[7423] = in[615] ^ in[222]; 
    assign layer_0[7424] = ~in[643]; 
    assign layer_0[7425] = ~(in[744] ^ in[481]); 
    assign layer_0[7426] = ~in[163] | (in[826] & in[163]); 
    assign layer_0[7427] = ~(in[603] ^ in[963]); 
    assign layer_0[7428] = in[730] | in[837]; 
    assign layer_0[7429] = in[85]; 
    assign layer_0[7430] = in[806] ^ in[731]; 
    assign layer_0[7431] = in[396] & in[375]; 
    assign layer_0[7432] = ~(in[743] ^ in[950]); 
    assign layer_0[7433] = in[822] ^ in[840]; 
    assign layer_0[7434] = 1'b1; 
    assign layer_0[7435] = in[604]; 
    assign layer_0[7436] = ~(in[935] ^ in[207]); 
    assign layer_0[7437] = in[582] ^ in[191]; 
    assign layer_0[7438] = ~in[854]; 
    assign layer_0[7439] = 1'b1; 
    assign layer_0[7440] = in[352] & ~in[629]; 
    assign layer_0[7441] = ~in[770]; 
    assign layer_0[7442] = in[1015] | in[500]; 
    assign layer_0[7443] = ~(in[835] ^ in[982]); 
    assign layer_0[7444] = ~in[617]; 
    assign layer_0[7445] = in[89] & in[228]; 
    assign layer_0[7446] = ~in[77] | (in[77] & in[504]); 
    assign layer_0[7447] = ~(in[790] ^ in[731]); 
    assign layer_0[7448] = ~(in[492] ^ in[905]); 
    assign layer_0[7449] = ~(in[235] ^ in[507]); 
    assign layer_0[7450] = ~in[622]; 
    assign layer_0[7451] = in[110] & in[502]; 
    assign layer_0[7452] = ~(in[972] & in[212]); 
    assign layer_0[7453] = in[609] | in[580]; 
    assign layer_0[7454] = in[185] & ~in[291]; 
    assign layer_0[7455] = ~(in[698] ^ in[963]); 
    assign layer_0[7456] = ~(in[156] ^ in[882]); 
    assign layer_0[7457] = in[518] & in[579]; 
    assign layer_0[7458] = in[1012] ^ in[627]; 
    assign layer_0[7459] = ~in[642] | (in[388] & in[642]); 
    assign layer_0[7460] = ~(in[148] & in[744]); 
    assign layer_0[7461] = in[122] ^ in[254]; 
    assign layer_0[7462] = ~in[744] | (in[252] & in[744]); 
    assign layer_0[7463] = in[476] & in[463]; 
    assign layer_0[7464] = ~in[78] | (in[78] & in[281]); 
    assign layer_0[7465] = ~(in[883] ^ in[508]); 
    assign layer_0[7466] = ~in[872] | (in[872] & in[880]); 
    assign layer_0[7467] = ~in[207] | (in[207] & in[685]); 
    assign layer_0[7468] = in[585] & ~in[1]; 
    assign layer_0[7469] = in[743] ^ in[853]; 
    assign layer_0[7470] = in[952] ^ in[548]; 
    assign layer_0[7471] = in[743] & ~in[595]; 
    assign layer_0[7472] = in[700] ^ in[501]; 
    assign layer_0[7473] = in[485] ^ in[840]; 
    assign layer_0[7474] = in[82]; 
    assign layer_0[7475] = ~in[870]; 
    assign layer_0[7476] = ~(in[522] ^ in[907]); 
    assign layer_0[7477] = in[60] & in[760]; 
    assign layer_0[7478] = ~in[70] | (in[257] & in[70]); 
    assign layer_0[7479] = ~in[380]; 
    assign layer_0[7480] = ~in[538]; 
    assign layer_0[7481] = ~(in[905] | in[747]); 
    assign layer_0[7482] = ~in[555]; 
    assign layer_0[7483] = in[741] | in[845]; 
    assign layer_0[7484] = in[193] ^ in[74]; 
    assign layer_0[7485] = in[301] ^ in[451]; 
    assign layer_0[7486] = in[844]; 
    assign layer_0[7487] = ~(in[365] | in[920]); 
    assign layer_0[7488] = ~in[634]; 
    assign layer_0[7489] = ~(in[788] ^ in[949]); 
    assign layer_0[7490] = ~(in[778] | in[458]); 
    assign layer_0[7491] = in[187] & in[103]; 
    assign layer_0[7492] = in[373] & in[452]; 
    assign layer_0[7493] = ~(in[659] ^ in[296]); 
    assign layer_0[7494] = ~in[581] | (in[581] & in[958]); 
    assign layer_0[7495] = ~(in[339] ^ in[873]); 
    assign layer_0[7496] = in[8]; 
    assign layer_0[7497] = in[317] ^ in[507]; 
    assign layer_0[7498] = in[788] & ~in[364]; 
    assign layer_0[7499] = in[821] | in[654]; 
    assign layer_0[7500] = in[601]; 
    assign layer_0[7501] = in[314] & in[583]; 
    assign layer_0[7502] = in[906] & ~in[731]; 
    assign layer_0[7503] = ~(in[824] & in[841]); 
    assign layer_0[7504] = ~(in[446] & in[512]); 
    assign layer_0[7505] = ~(in[765] | in[540]); 
    assign layer_0[7506] = in[276] & ~in[961]; 
    assign layer_0[7507] = ~(in[601] ^ in[799]); 
    assign layer_0[7508] = in[452] & ~in[621]; 
    assign layer_0[7509] = ~in[655] | (in[611] & in[655]); 
    assign layer_0[7510] = ~(in[617] ^ in[791]); 
    assign layer_0[7511] = in[659] | in[49]; 
    assign layer_0[7512] = ~(in[100] ^ in[612]); 
    assign layer_0[7513] = ~in[875] | (in[30] & in[875]); 
    assign layer_0[7514] = ~(in[368] | in[525]); 
    assign layer_0[7515] = ~(in[117] & in[216]); 
    assign layer_0[7516] = ~(in[646] ^ in[7]); 
    assign layer_0[7517] = ~(in[806] ^ in[261]); 
    assign layer_0[7518] = in[112] ^ in[218]; 
    assign layer_0[7519] = ~in[725] | (in[597] & in[725]); 
    assign layer_0[7520] = ~(in[835] ^ in[773]); 
    assign layer_0[7521] = in[591] ^ in[699]; 
    assign layer_0[7522] = in[766] ^ in[873]; 
    assign layer_0[7523] = ~(in[974] | in[247]); 
    assign layer_0[7524] = in[135] & ~in[628]; 
    assign layer_0[7525] = ~(in[275] ^ in[350]); 
    assign layer_0[7526] = 1'b0; 
    assign layer_0[7527] = ~(in[775] | in[648]); 
    assign layer_0[7528] = in[820] & ~in[212]; 
    assign layer_0[7529] = ~(in[953] | in[713]); 
    assign layer_0[7530] = in[308] & ~in[510]; 
    assign layer_0[7531] = ~(in[615] & in[649]); 
    assign layer_0[7532] = in[92] & ~in[643]; 
    assign layer_0[7533] = ~(in[828] ^ in[387]); 
    assign layer_0[7534] = in[904] & ~in[273]; 
    assign layer_0[7535] = ~in[308] | (in[10] & in[308]); 
    assign layer_0[7536] = in[575] ^ in[415]; 
    assign layer_0[7537] = ~(in[902] | in[477]); 
    assign layer_0[7538] = in[962] & in[883]; 
    assign layer_0[7539] = in[51] & in[939]; 
    assign layer_0[7540] = ~in[46] | (in[637] & in[46]); 
    assign layer_0[7541] = in[825] & ~in[577]; 
    assign layer_0[7542] = in[455] & in[1018]; 
    assign layer_0[7543] = ~(in[665] & in[444]); 
    assign layer_0[7544] = ~in[303]; 
    assign layer_0[7545] = in[890] & ~in[795]; 
    assign layer_0[7546] = ~(in[663] & in[260]); 
    assign layer_0[7547] = in[749] & ~in[907]; 
    assign layer_0[7548] = ~in[522] | (in[956] & in[522]); 
    assign layer_0[7549] = ~in[521]; 
    assign layer_0[7550] = in[887]; 
    assign layer_0[7551] = in[909] & ~in[751]; 
    assign layer_0[7552] = in[922] ^ in[842]; 
    assign layer_0[7553] = ~(in[315] & in[984]); 
    assign layer_0[7554] = ~(in[19] | in[571]); 
    assign layer_0[7555] = in[628] & ~in[860]; 
    assign layer_0[7556] = in[685] & ~in[359]; 
    assign layer_0[7557] = ~(in[866] ^ in[840]); 
    assign layer_0[7558] = ~in[168] | (in[654] & in[168]); 
    assign layer_0[7559] = in[540]; 
    assign layer_0[7560] = in[634] & in[714]; 
    assign layer_0[7561] = ~in[610]; 
    assign layer_0[7562] = in[324]; 
    assign layer_0[7563] = ~in[520]; 
    assign layer_0[7564] = ~in[828]; 
    assign layer_0[7565] = in[440]; 
    assign layer_0[7566] = ~(in[956] ^ in[469]); 
    assign layer_0[7567] = ~in[475] | (in[723] & in[475]); 
    assign layer_0[7568] = in[899] ^ in[900]; 
    assign layer_0[7569] = ~(in[210] ^ in[300]); 
    assign layer_0[7570] = in[936] ^ in[901]; 
    assign layer_0[7571] = in[969] & ~in[349]; 
    assign layer_0[7572] = ~(in[517] ^ in[291]); 
    assign layer_0[7573] = in[890] ^ in[76]; 
    assign layer_0[7574] = in[876] ^ in[843]; 
    assign layer_0[7575] = ~(in[1000] ^ in[1002]); 
    assign layer_0[7576] = ~in[49]; 
    assign layer_0[7577] = in[41]; 
    assign layer_0[7578] = ~in[794] | (in[1003] & in[794]); 
    assign layer_0[7579] = ~(in[817] & in[774]); 
    assign layer_0[7580] = in[293] & in[488]; 
    assign layer_0[7581] = in[713]; 
    assign layer_0[7582] = ~(in[12] ^ in[674]); 
    assign layer_0[7583] = in[827] ^ in[722]; 
    assign layer_0[7584] = in[482]; 
    assign layer_0[7585] = ~(in[967] ^ in[939]); 
    assign layer_0[7586] = ~in[46] | (in[46] & in[239]); 
    assign layer_0[7587] = ~in[474]; 
    assign layer_0[7588] = ~(in[981] ^ in[207]); 
    assign layer_0[7589] = in[428] ^ in[66]; 
    assign layer_0[7590] = in[898] & in[974]; 
    assign layer_0[7591] = in[584] & in[427]; 
    assign layer_0[7592] = in[931]; 
    assign layer_0[7593] = in[230] & ~in[705]; 
    assign layer_0[7594] = ~(in[95] | in[532]); 
    assign layer_0[7595] = ~in[842]; 
    assign layer_0[7596] = in[432]; 
    assign layer_0[7597] = in[760] ^ in[613]; 
    assign layer_0[7598] = ~in[500] | (in[956] & in[500]); 
    assign layer_0[7599] = ~in[260] | (in[830] & in[260]); 
    assign layer_0[7600] = in[84]; 
    assign layer_0[7601] = in[140] & ~in[303]; 
    assign layer_0[7602] = ~(in[92] ^ in[518]); 
    assign layer_0[7603] = in[45] ^ in[549]; 
    assign layer_0[7604] = ~(in[534] ^ in[242]); 
    assign layer_0[7605] = ~in[806] | (in[79] & in[806]); 
    assign layer_0[7606] = 1'b0; 
    assign layer_0[7607] = ~in[708] | (in[930] & in[708]); 
    assign layer_0[7608] = ~(in[673] & in[191]); 
    assign layer_0[7609] = ~(in[356] ^ in[788]); 
    assign layer_0[7610] = ~(in[358] ^ in[627]); 
    assign layer_0[7611] = in[843] & in[623]; 
    assign layer_0[7612] = in[412] & in[1016]; 
    assign layer_0[7613] = ~(in[885] ^ in[760]); 
    assign layer_0[7614] = ~(in[210] & in[967]); 
    assign layer_0[7615] = in[314]; 
    assign layer_0[7616] = in[841] ^ in[750]; 
    assign layer_0[7617] = in[276] ^ in[435]; 
    assign layer_0[7618] = ~in[620]; 
    assign layer_0[7619] = ~in[535]; 
    assign layer_0[7620] = ~in[627] | (in[259] & in[627]); 
    assign layer_0[7621] = in[860] ^ in[995]; 
    assign layer_0[7622] = in[916] | in[999]; 
    assign layer_0[7623] = in[635] & ~in[731]; 
    assign layer_0[7624] = in[401] & in[926]; 
    assign layer_0[7625] = in[634] & in[621]; 
    assign layer_0[7626] = in[531]; 
    assign layer_0[7627] = ~(in[50] ^ in[836]); 
    assign layer_0[7628] = ~(in[774] | in[792]); 
    assign layer_0[7629] = in[518] & ~in[651]; 
    assign layer_0[7630] = ~(in[341] | in[676]); 
    assign layer_0[7631] = ~in[491] | (in[491] & in[1014]); 
    assign layer_0[7632] = ~(in[627] ^ in[414]); 
    assign layer_0[7633] = in[633] ^ in[613]; 
    assign layer_0[7634] = ~(in[838] ^ in[810]); 
    assign layer_0[7635] = in[518] ^ in[946]; 
    assign layer_0[7636] = in[905]; 
    assign layer_0[7637] = ~(in[48] ^ in[473]); 
    assign layer_0[7638] = in[378] ^ in[757]; 
    assign layer_0[7639] = ~(in[30] | in[796]); 
    assign layer_0[7640] = 1'b0; 
    assign layer_0[7641] = ~(in[902] ^ in[917]); 
    assign layer_0[7642] = ~in[488]; 
    assign layer_0[7643] = ~(in[856] & in[940]); 
    assign layer_0[7644] = ~in[520] | (in[13] & in[520]); 
    assign layer_0[7645] = in[903] ^ in[653]; 
    assign layer_0[7646] = in[673] ^ in[726]; 
    assign layer_0[7647] = ~(in[264] ^ in[94]); 
    assign layer_0[7648] = in[649] ^ in[732]; 
    assign layer_0[7649] = in[170] & ~in[826]; 
    assign layer_0[7650] = in[193]; 
    assign layer_0[7651] = ~(in[881] & in[721]); 
    assign layer_0[7652] = ~(in[366] ^ in[455]); 
    assign layer_0[7653] = ~(in[317] | in[256]); 
    assign layer_0[7654] = ~in[50]; 
    assign layer_0[7655] = in[724] ^ in[948]; 
    assign layer_0[7656] = ~in[216] | (in[222] & in[216]); 
    assign layer_0[7657] = in[655]; 
    assign layer_0[7658] = ~in[407]; 
    assign layer_0[7659] = ~(in[400] | in[727]); 
    assign layer_0[7660] = ~(in[547] ^ in[365]); 
    assign layer_0[7661] = ~(in[571] ^ in[739]); 
    assign layer_0[7662] = in[569] & ~in[809]; 
    assign layer_0[7663] = ~(in[318] ^ in[842]); 
    assign layer_0[7664] = ~(in[757] | in[794]); 
    assign layer_0[7665] = ~in[597] | (in[972] & in[597]); 
    assign layer_0[7666] = in[8]; 
    assign layer_0[7667] = ~(in[885] ^ in[980]); 
    assign layer_0[7668] = ~(in[681] ^ in[808]); 
    assign layer_0[7669] = in[739] ^ in[548]; 
    assign layer_0[7670] = ~(in[910] ^ in[216]); 
    assign layer_0[7671] = in[696] ^ in[888]; 
    assign layer_0[7672] = in[370] ^ in[465]; 
    assign layer_0[7673] = ~in[825]; 
    assign layer_0[7674] = ~(in[163] & in[54]); 
    assign layer_0[7675] = ~(in[199] & in[303]); 
    assign layer_0[7676] = ~(in[419] ^ in[175]); 
    assign layer_0[7677] = 1'b1; 
    assign layer_0[7678] = in[836] ^ in[663]; 
    assign layer_0[7679] = ~in[274] | (in[274] & in[796]); 
    assign layer_0[7680] = in[654]; 
    assign layer_0[7681] = ~(in[193] | in[747]); 
    assign layer_0[7682] = in[573] | in[981]; 
    assign layer_0[7683] = in[840] ^ in[730]; 
    assign layer_0[7684] = ~in[859] | (in[649] & in[859]); 
    assign layer_0[7685] = in[821] | in[824]; 
    assign layer_0[7686] = ~in[34]; 
    assign layer_0[7687] = in[541] & in[199]; 
    assign layer_0[7688] = ~(in[999] | in[323]); 
    assign layer_0[7689] = 1'b1; 
    assign layer_0[7690] = in[487] & ~in[96]; 
    assign layer_0[7691] = in[1009] ^ in[380]; 
    assign layer_0[7692] = ~(in[451] ^ in[51]); 
    assign layer_0[7693] = in[588] | in[953]; 
    assign layer_0[7694] = ~(in[1000] ^ in[493]); 
    assign layer_0[7695] = in[711] ^ in[557]; 
    assign layer_0[7696] = in[33] | in[874]; 
    assign layer_0[7697] = in[119] & ~in[821]; 
    assign layer_0[7698] = in[417] & ~in[41]; 
    assign layer_0[7699] = in[724] ^ in[844]; 
    assign layer_0[7700] = in[125] & in[922]; 
    assign layer_0[7701] = in[672] ^ in[40]; 
    assign layer_0[7702] = ~(in[396] ^ in[158]); 
    assign layer_0[7703] = in[310]; 
    assign layer_0[7704] = in[398] ^ in[242]; 
    assign layer_0[7705] = in[548] & ~in[707]; 
    assign layer_0[7706] = ~in[990]; 
    assign layer_0[7707] = ~(in[477] ^ in[652]); 
    assign layer_0[7708] = in[679] & ~in[568]; 
    assign layer_0[7709] = in[620] ^ in[267]; 
    assign layer_0[7710] = ~(in[655] ^ in[474]); 
    assign layer_0[7711] = ~in[450]; 
    assign layer_0[7712] = ~in[938] | (in[938] & in[96]); 
    assign layer_0[7713] = in[18] ^ in[758]; 
    assign layer_0[7714] = in[707] ^ in[587]; 
    assign layer_0[7715] = in[582] ^ in[554]; 
    assign layer_0[7716] = ~(in[502] | in[978]); 
    assign layer_0[7717] = ~in[259] | (in[555] & in[259]); 
    assign layer_0[7718] = ~(in[620] | in[1000]); 
    assign layer_0[7719] = in[901] | in[900]; 
    assign layer_0[7720] = ~(in[743] & in[510]); 
    assign layer_0[7721] = in[142] ^ in[69]; 
    assign layer_0[7722] = ~in[552]; 
    assign layer_0[7723] = ~(in[643] ^ in[158]); 
    assign layer_0[7724] = ~(in[363] ^ in[689]); 
    assign layer_0[7725] = ~in[957] | (in[522] & in[957]); 
    assign layer_0[7726] = in[387] | in[913]; 
    assign layer_0[7727] = in[579]; 
    assign layer_0[7728] = ~in[691]; 
    assign layer_0[7729] = ~(in[676] ^ in[157]); 
    assign layer_0[7730] = in[875]; 
    assign layer_0[7731] = ~(in[493] & in[723]); 
    assign layer_0[7732] = ~in[458] | (in[614] & in[458]); 
    assign layer_0[7733] = 1'b1; 
    assign layer_0[7734] = ~(in[384] ^ in[726]); 
    assign layer_0[7735] = ~(in[941] ^ in[590]); 
    assign layer_0[7736] = ~in[648] | (in[648] & in[613]); 
    assign layer_0[7737] = ~(in[141] & in[603]); 
    assign layer_0[7738] = in[164] & ~in[139]; 
    assign layer_0[7739] = in[583] ^ in[905]; 
    assign layer_0[7740] = ~(in[972] ^ in[209]); 
    assign layer_0[7741] = in[746] & ~in[354]; 
    assign layer_0[7742] = in[413] ^ in[315]; 
    assign layer_0[7743] = in[903] & in[217]; 
    assign layer_0[7744] = ~in[388]; 
    assign layer_0[7745] = ~in[288]; 
    assign layer_0[7746] = ~(in[914] ^ in[763]); 
    assign layer_0[7747] = ~(in[615] ^ in[102]); 
    assign layer_0[7748] = ~in[442] | (in[920] & in[442]); 
    assign layer_0[7749] = in[615] ^ in[427]; 
    assign layer_0[7750] = ~in[297]; 
    assign layer_0[7751] = ~in[496]; 
    assign layer_0[7752] = ~(in[825] & in[889]); 
    assign layer_0[7753] = ~in[825] | (in[825] & in[805]); 
    assign layer_0[7754] = in[504]; 
    assign layer_0[7755] = in[746] ^ in[81]; 
    assign layer_0[7756] = ~(in[839] ^ in[486]); 
    assign layer_0[7757] = in[597] | in[459]; 
    assign layer_0[7758] = ~(in[948] ^ in[941]); 
    assign layer_0[7759] = in[367] ^ in[686]; 
    assign layer_0[7760] = ~(in[1020] ^ in[939]); 
    assign layer_0[7761] = in[346] & ~in[596]; 
    assign layer_0[7762] = ~in[316] | (in[790] & in[316]); 
    assign layer_0[7763] = ~in[536]; 
    assign layer_0[7764] = ~(in[638] & in[662]); 
    assign layer_0[7765] = ~in[567] | (in[567] & in[741]); 
    assign layer_0[7766] = in[638] & ~in[418]; 
    assign layer_0[7767] = in[904] ^ in[243]; 
    assign layer_0[7768] = in[596] ^ in[636]; 
    assign layer_0[7769] = in[51]; 
    assign layer_0[7770] = in[908] & ~in[902]; 
    assign layer_0[7771] = ~in[641]; 
    assign layer_0[7772] = in[111] & ~in[510]; 
    assign layer_0[7773] = in[357]; 
    assign layer_0[7774] = in[4] & in[723]; 
    assign layer_0[7775] = ~(in[571] ^ in[112]); 
    assign layer_0[7776] = ~(in[501] ^ in[916]); 
    assign layer_0[7777] = in[567] & ~in[124]; 
    assign layer_0[7778] = in[902]; 
    assign layer_0[7779] = in[381] ^ in[729]; 
    assign layer_0[7780] = ~in[792] | (in[80] & in[792]); 
    assign layer_0[7781] = in[810] | in[572]; 
    assign layer_0[7782] = ~(in[938] ^ in[614]); 
    assign layer_0[7783] = in[307] & in[259]; 
    assign layer_0[7784] = in[856] | in[668]; 
    assign layer_0[7785] = in[561]; 
    assign layer_0[7786] = ~(in[97] ^ in[84]); 
    assign layer_0[7787] = in[839] ^ in[654]; 
    assign layer_0[7788] = ~in[119] | (in[747] & in[119]); 
    assign layer_0[7789] = ~(in[933] ^ in[537]); 
    assign layer_0[7790] = in[34] & ~in[702]; 
    assign layer_0[7791] = ~(in[507] ^ in[619]); 
    assign layer_0[7792] = in[611] ^ in[337]; 
    assign layer_0[7793] = ~(in[142] ^ in[197]); 
    assign layer_0[7794] = in[642] ^ in[895]; 
    assign layer_0[7795] = ~in[852] | (in[592] & in[852]); 
    assign layer_0[7796] = in[629] ^ in[756]; 
    assign layer_0[7797] = ~(in[356] & in[457]); 
    assign layer_0[7798] = in[689] | in[759]; 
    assign layer_0[7799] = in[950] & ~in[210]; 
    assign layer_0[7800] = in[853] | in[142]; 
    assign layer_0[7801] = in[63] & ~in[943]; 
    assign layer_0[7802] = ~(in[372] ^ in[634]); 
    assign layer_0[7803] = in[578] | in[460]; 
    assign layer_0[7804] = ~in[459] | (in[611] & in[459]); 
    assign layer_0[7805] = ~(in[707] ^ in[323]); 
    assign layer_0[7806] = in[73] ^ in[604]; 
    assign layer_0[7807] = ~in[23] | (in[23] & in[909]); 
    assign layer_0[7808] = in[933]; 
    assign layer_0[7809] = ~(in[1017] ^ in[663]); 
    assign layer_0[7810] = in[578] | in[712]; 
    assign layer_0[7811] = in[934] ^ in[311]; 
    assign layer_0[7812] = in[938] | in[613]; 
    assign layer_0[7813] = in[808]; 
    assign layer_0[7814] = in[374] & ~in[12]; 
    assign layer_0[7815] = ~in[410] | (in[5] & in[410]); 
    assign layer_0[7816] = in[3] & ~in[957]; 
    assign layer_0[7817] = in[857] & ~in[817]; 
    assign layer_0[7818] = ~(in[344] ^ in[502]); 
    assign layer_0[7819] = ~(in[631] ^ in[699]); 
    assign layer_0[7820] = in[745] & ~in[892]; 
    assign layer_0[7821] = ~in[595]; 
    assign layer_0[7822] = ~(in[949] ^ in[715]); 
    assign layer_0[7823] = in[354] & ~in[318]; 
    assign layer_0[7824] = ~(in[699] ^ in[280]); 
    assign layer_0[7825] = 1'b1; 
    assign layer_0[7826] = ~in[581]; 
    assign layer_0[7827] = ~(in[621] ^ in[712]); 
    assign layer_0[7828] = ~in[875]; 
    assign layer_0[7829] = ~(in[263] | in[965]); 
    assign layer_0[7830] = in[953]; 
    assign layer_0[7831] = ~in[864] | (in[864] & in[752]); 
    assign layer_0[7832] = ~(in[188] | in[1000]); 
    assign layer_0[7833] = ~(in[762] & in[118]); 
    assign layer_0[7834] = in[970] & ~in[264]; 
    assign layer_0[7835] = ~in[867]; 
    assign layer_0[7836] = in[448] ^ in[886]; 
    assign layer_0[7837] = ~(in[109] ^ in[419]); 
    assign layer_0[7838] = ~(in[105] & in[636]); 
    assign layer_0[7839] = ~(in[580] ^ in[582]); 
    assign layer_0[7840] = ~in[640]; 
    assign layer_0[7841] = in[757]; 
    assign layer_0[7842] = in[996]; 
    assign layer_0[7843] = ~in[634] | (in[634] & in[596]); 
    assign layer_0[7844] = in[819] | in[654]; 
    assign layer_0[7845] = ~(in[536] ^ in[843]); 
    assign layer_0[7846] = in[661] & in[226]; 
    assign layer_0[7847] = ~(in[61] ^ in[460]); 
    assign layer_0[7848] = ~in[739]; 
    assign layer_0[7849] = in[364] & in[149]; 
    assign layer_0[7850] = ~(in[974] & in[1002]); 
    assign layer_0[7851] = ~(in[457] & in[329]); 
    assign layer_0[7852] = ~(in[115] ^ in[347]); 
    assign layer_0[7853] = in[872]; 
    assign layer_0[7854] = in[651] & ~in[706]; 
    assign layer_0[7855] = ~in[99] | (in[79] & in[99]); 
    assign layer_0[7856] = in[968] ^ in[776]; 
    assign layer_0[7857] = in[115] & ~in[668]; 
    assign layer_0[7858] = in[263] ^ in[728]; 
    assign layer_0[7859] = in[778] ^ in[807]; 
    assign layer_0[7860] = in[485] | in[719]; 
    assign layer_0[7861] = in[918] ^ in[804]; 
    assign layer_0[7862] = ~(in[927] | in[964]); 
    assign layer_0[7863] = in[587] ^ in[790]; 
    assign layer_0[7864] = in[764] | in[698]; 
    assign layer_0[7865] = in[963] & ~in[304]; 
    assign layer_0[7866] = in[694] & ~in[774]; 
    assign layer_0[7867] = in[883] & in[238]; 
    assign layer_0[7868] = in[301]; 
    assign layer_0[7869] = in[744] & in[308]; 
    assign layer_0[7870] = in[954] | in[853]; 
    assign layer_0[7871] = in[22] & in[362]; 
    assign layer_0[7872] = 1'b1; 
    assign layer_0[7873] = in[709] ^ in[634]; 
    assign layer_0[7874] = in[298] & ~in[473]; 
    assign layer_0[7875] = ~in[634] | (in[634] & in[980]); 
    assign layer_0[7876] = ~in[660] | (in[870] & in[660]); 
    assign layer_0[7877] = in[971]; 
    assign layer_0[7878] = ~in[630]; 
    assign layer_0[7879] = ~(in[77] ^ in[254]); 
    assign layer_0[7880] = ~(in[612] ^ in[952]); 
    assign layer_0[7881] = in[611] & ~in[566]; 
    assign layer_0[7882] = ~in[253]; 
    assign layer_0[7883] = in[495] ^ in[1022]; 
    assign layer_0[7884] = ~(in[585] ^ in[1009]); 
    assign layer_0[7885] = ~in[371]; 
    assign layer_0[7886] = ~(in[699] | in[715]); 
    assign layer_0[7887] = ~in[416]; 
    assign layer_0[7888] = ~(in[547] | in[28]); 
    assign layer_0[7889] = in[1020] ^ in[140]; 
    assign layer_0[7890] = ~in[299]; 
    assign layer_0[7891] = in[2] | in[499]; 
    assign layer_0[7892] = ~in[875] | (in[875] & in[944]); 
    assign layer_0[7893] = ~in[733] | (in[573] & in[733]); 
    assign layer_0[7894] = ~(in[958] & in[934]); 
    assign layer_0[7895] = in[68]; 
    assign layer_0[7896] = in[503] ^ in[501]; 
    assign layer_0[7897] = in[247]; 
    assign layer_0[7898] = ~in[374]; 
    assign layer_0[7899] = in[71] & ~in[467]; 
    assign layer_0[7900] = in[76] & in[299]; 
    assign layer_0[7901] = ~in[979] | (in[979] & in[18]); 
    assign layer_0[7902] = ~in[19]; 
    assign layer_0[7903] = in[684] & ~in[264]; 
    assign layer_0[7904] = ~in[886] | (in[788] & in[886]); 
    assign layer_0[7905] = in[810] ^ in[614]; 
    assign layer_0[7906] = in[231]; 
    assign layer_0[7907] = in[603] & ~in[612]; 
    assign layer_0[7908] = ~(in[697] ^ in[649]); 
    assign layer_0[7909] = ~(in[612] ^ in[604]); 
    assign layer_0[7910] = ~(in[492] ^ in[842]); 
    assign layer_0[7911] = in[1021] ^ in[30]; 
    assign layer_0[7912] = ~(in[17] & in[775]); 
    assign layer_0[7913] = ~(in[264] | in[264]); 
    assign layer_0[7914] = in[3] ^ in[136]; 
    assign layer_0[7915] = in[702] ^ in[582]; 
    assign layer_0[7916] = ~(in[301] | in[506]); 
    assign layer_0[7917] = in[420] & ~in[19]; 
    assign layer_0[7918] = ~(in[744] ^ in[923]); 
    assign layer_0[7919] = ~in[659] | (in[659] & in[680]); 
    assign layer_0[7920] = ~(in[937] ^ in[999]); 
    assign layer_0[7921] = ~in[504] | (in[565] & in[504]); 
    assign layer_0[7922] = ~in[391]; 
    assign layer_0[7923] = ~(in[789] ^ in[535]); 
    assign layer_0[7924] = ~(in[882] | in[280]); 
    assign layer_0[7925] = in[821] | in[312]; 
    assign layer_0[7926] = ~(in[556] ^ in[534]); 
    assign layer_0[7927] = ~in[493] | (in[476] & in[493]); 
    assign layer_0[7928] = in[540] ^ in[521]; 
    assign layer_0[7929] = ~(in[819] ^ in[862]); 
    assign layer_0[7930] = ~(in[419] & in[614]); 
    assign layer_0[7931] = ~(in[658] ^ in[211]); 
    assign layer_0[7932] = ~in[965] | (in[34] & in[965]); 
    assign layer_0[7933] = in[632] & in[687]; 
    assign layer_0[7934] = in[608] | in[952]; 
    assign layer_0[7935] = in[252]; 
    assign layer_0[7936] = in[465] & in[894]; 
    assign layer_0[7937] = ~in[805] | (in[805] & in[556]); 
    assign layer_0[7938] = in[892]; 
    assign layer_0[7939] = ~(in[655] | in[404]); 
    assign layer_0[7940] = in[751] | in[229]; 
    assign layer_0[7941] = in[725] ^ in[483]; 
    assign layer_0[7942] = ~(in[66] ^ in[858]); 
    assign layer_0[7943] = in[752] | in[760]; 
    assign layer_0[7944] = in[21] & ~in[950]; 
    assign layer_0[7945] = ~(in[30] ^ in[264]); 
    assign layer_0[7946] = ~(in[889] ^ in[918]); 
    assign layer_0[7947] = ~(in[1016] ^ in[176]); 
    assign layer_0[7948] = ~(in[473] ^ in[715]); 
    assign layer_0[7949] = in[252] & ~in[865]; 
    assign layer_0[7950] = in[508] ^ in[876]; 
    assign layer_0[7951] = ~(in[448] | in[629]); 
    assign layer_0[7952] = ~(in[74] & in[450]); 
    assign layer_0[7953] = ~(in[890] & in[825]); 
    assign layer_0[7954] = in[239] & ~in[1004]; 
    assign layer_0[7955] = in[156] & ~in[740]; 
    assign layer_0[7956] = in[276] ^ in[548]; 
    assign layer_0[7957] = in[934] ^ in[4]; 
    assign layer_0[7958] = ~in[132]; 
    assign layer_0[7959] = in[505] | in[888]; 
    assign layer_0[7960] = ~in[403] | (in[403] & in[676]); 
    assign layer_0[7961] = ~in[541] | (in[1006] & in[541]); 
    assign layer_0[7962] = in[92] ^ in[268]; 
    assign layer_0[7963] = ~(in[930] ^ in[316]); 
    assign layer_0[7964] = in[670] & ~in[804]; 
    assign layer_0[7965] = ~in[404] | (in[404] & in[210]); 
    assign layer_0[7966] = ~(in[223] ^ in[404]); 
    assign layer_0[7967] = in[219] & ~in[891]; 
    assign layer_0[7968] = in[315] ^ in[687]; 
    assign layer_0[7969] = in[96] | in[845]; 
    assign layer_0[7970] = in[627]; 
    assign layer_0[7971] = in[451] | in[939]; 
    assign layer_0[7972] = in[733] ^ in[961]; 
    assign layer_0[7973] = in[873] ^ in[759]; 
    assign layer_0[7974] = in[903] & ~in[651]; 
    assign layer_0[7975] = in[349] ^ in[1012]; 
    assign layer_0[7976] = in[563]; 
    assign layer_0[7977] = ~in[833]; 
    assign layer_0[7978] = in[403]; 
    assign layer_0[7979] = in[84] | in[293]; 
    assign layer_0[7980] = ~in[440] | (in[440] & in[998]); 
    assign layer_0[7981] = in[731] ^ in[175]; 
    assign layer_0[7982] = ~in[735]; 
    assign layer_0[7983] = ~(in[314] & in[487]); 
    assign layer_0[7984] = in[1016] | in[812]; 
    assign layer_0[7985] = in[955] & ~in[253]; 
    assign layer_0[7986] = in[598] ^ in[596]; 
    assign layer_0[7987] = ~(in[596] ^ in[284]); 
    assign layer_0[7988] = ~(in[641] ^ in[777]); 
    assign layer_0[7989] = ~in[348] | (in[356] & in[348]); 
    assign layer_0[7990] = in[446] & ~in[878]; 
    assign layer_0[7991] = ~(in[33] ^ in[308]); 
    assign layer_0[7992] = in[40] | in[34]; 
    assign layer_0[7993] = ~(in[371] ^ in[870]); 
    assign layer_0[7994] = in[411] & ~in[552]; 
    assign layer_0[7995] = in[466] & in[310]; 
    assign layer_0[7996] = ~(in[600] ^ in[599]); 
    assign layer_0[7997] = in[660] | in[915]; 
    assign layer_0[7998] = in[938] | in[238]; 
    assign layer_0[7999] = in[122] & ~in[792]; 
    assign layer_0[8000] = in[874] | in[732]; 
    assign layer_0[8001] = ~(in[915] ^ in[551]); 
    assign layer_0[8002] = ~in[900]; 
    assign layer_0[8003] = ~(in[596] | in[619]); 
    assign layer_0[8004] = ~(in[656] ^ in[649]); 
    assign layer_0[8005] = in[974] ^ in[117]; 
    assign layer_0[8006] = ~(in[934] ^ in[919]); 
    assign layer_0[8007] = ~(in[446] ^ in[293]); 
    assign layer_0[8008] = in[243] ^ in[606]; 
    assign layer_0[8009] = in[445] & in[984]; 
    assign layer_0[8010] = ~in[731]; 
    assign layer_0[8011] = in[863] ^ in[856]; 
    assign layer_0[8012] = ~in[1002] | (in[451] & in[1002]); 
    assign layer_0[8013] = in[264] & ~in[403]; 
    assign layer_0[8014] = ~(in[667] ^ in[731]); 
    assign layer_0[8015] = in[633] & ~in[502]; 
    assign layer_0[8016] = ~(in[724] ^ in[390]); 
    assign layer_0[8017] = in[498]; 
    assign layer_0[8018] = ~(in[41] & in[755]); 
    assign layer_0[8019] = in[6] & ~in[126]; 
    assign layer_0[8020] = ~in[835] | (in[835] & in[968]); 
    assign layer_0[8021] = ~(in[508] ^ in[919]); 
    assign layer_0[8022] = ~(in[607] & in[408]); 
    assign layer_0[8023] = in[267]; 
    assign layer_0[8024] = ~(in[478] & in[1016]); 
    assign layer_0[8025] = in[629] ^ in[101]; 
    assign layer_0[8026] = in[344] & ~in[898]; 
    assign layer_0[8027] = in[894] & in[489]; 
    assign layer_0[8028] = ~(in[21] | in[175]); 
    assign layer_0[8029] = ~in[163]; 
    assign layer_0[8030] = in[449]; 
    assign layer_0[8031] = in[63] & ~in[754]; 
    assign layer_0[8032] = ~(in[609] | in[667]); 
    assign layer_0[8033] = ~(in[886] ^ in[869]); 
    assign layer_0[8034] = ~(in[18] ^ in[631]); 
    assign layer_0[8035] = ~in[701] | (in[701] & in[69]); 
    assign layer_0[8036] = ~(in[567] ^ in[813]); 
    assign layer_0[8037] = in[535] & ~in[633]; 
    assign layer_0[8038] = ~in[795]; 
    assign layer_0[8039] = in[3] ^ in[823]; 
    assign layer_0[8040] = ~(in[888] | in[252]); 
    assign layer_0[8041] = ~in[28]; 
    assign layer_0[8042] = in[286]; 
    assign layer_0[8043] = in[97] & in[112]; 
    assign layer_0[8044] = ~in[661]; 
    assign layer_0[8045] = in[445] ^ in[434]; 
    assign layer_0[8046] = in[763] | in[316]; 
    assign layer_0[8047] = ~in[646] | (in[646] & in[572]); 
    assign layer_0[8048] = in[603]; 
    assign layer_0[8049] = ~(in[301] ^ in[20]); 
    assign layer_0[8050] = ~(in[819] ^ in[179]); 
    assign layer_0[8051] = in[678] & ~in[1017]; 
    assign layer_0[8052] = ~(in[758] ^ in[761]); 
    assign layer_0[8053] = in[797] | in[20]; 
    assign layer_0[8054] = ~(in[648] & in[638]); 
    assign layer_0[8055] = in[282] & in[266]; 
    assign layer_0[8056] = in[131]; 
    assign layer_0[8057] = in[428] & ~in[779]; 
    assign layer_0[8058] = ~(in[599] ^ in[823]); 
    assign layer_0[8059] = 1'b1; 
    assign layer_0[8060] = in[812] | in[470]; 
    assign layer_0[8061] = in[569] & ~in[844]; 
    assign layer_0[8062] = in[924] ^ in[522]; 
    assign layer_0[8063] = in[100] | in[867]; 
    assign layer_0[8064] = ~(in[111] ^ in[275]); 
    assign layer_0[8065] = ~(in[869] ^ in[386]); 
    assign layer_0[8066] = ~in[305] | (in[305] & in[1009]); 
    assign layer_0[8067] = in[338]; 
    assign layer_0[8068] = in[804]; 
    assign layer_0[8069] = ~(in[548] | in[900]); 
    assign layer_0[8070] = in[487] ^ in[710]; 
    assign layer_0[8071] = ~(in[707] ^ in[904]); 
    assign layer_0[8072] = in[409] & ~in[986]; 
    assign layer_0[8073] = ~(in[743] ^ in[368]); 
    assign layer_0[8074] = in[531] | in[630]; 
    assign layer_0[8075] = in[395] & ~in[36]; 
    assign layer_0[8076] = ~(in[612] ^ in[980]); 
    assign layer_0[8077] = ~(in[855] & in[365]); 
    assign layer_0[8078] = ~(in[91] & in[825]); 
    assign layer_0[8079] = ~in[572]; 
    assign layer_0[8080] = in[857] & ~in[966]; 
    assign layer_0[8081] = ~(in[493] ^ in[207]); 
    assign layer_0[8082] = in[819] | in[465]; 
    assign layer_0[8083] = in[876]; 
    assign layer_0[8084] = in[925] ^ in[232]; 
    assign layer_0[8085] = ~in[368]; 
    assign layer_0[8086] = in[101] ^ in[703]; 
    assign layer_0[8087] = ~(in[664] & in[228]); 
    assign layer_0[8088] = in[618] ^ in[855]; 
    assign layer_0[8089] = ~in[754]; 
    assign layer_0[8090] = in[49]; 
    assign layer_0[8091] = ~in[556] | (in[700] & in[556]); 
    assign layer_0[8092] = ~in[858] | (in[178] & in[858]); 
    assign layer_0[8093] = ~in[356] | (in[356] & in[986]); 
    assign layer_0[8094] = in[723] & ~in[677]; 
    assign layer_0[8095] = ~(in[489] ^ in[789]); 
    assign layer_0[8096] = in[613] & ~in[611]; 
    assign layer_0[8097] = ~in[111]; 
    assign layer_0[8098] = ~(in[858] ^ in[837]); 
    assign layer_0[8099] = ~(in[706] ^ in[629]); 
    assign layer_0[8100] = in[753] ^ in[283]; 
    assign layer_0[8101] = ~(in[730] & in[726]); 
    assign layer_0[8102] = ~(in[740] & in[406]); 
    assign layer_0[8103] = ~(in[937] ^ in[938]); 
    assign layer_0[8104] = ~(in[967] ^ in[568]); 
    assign layer_0[8105] = ~(in[612] ^ in[603]); 
    assign layer_0[8106] = ~in[82]; 
    assign layer_0[8107] = in[806] ^ in[660]; 
    assign layer_0[8108] = in[596]; 
    assign layer_0[8109] = ~(in[701] | in[926]); 
    assign layer_0[8110] = in[588] ^ in[508]; 
    assign layer_0[8111] = ~in[775] | (in[775] & in[820]); 
    assign layer_0[8112] = ~in[1016]; 
    assign layer_0[8113] = ~(in[973] ^ in[870]); 
    assign layer_0[8114] = ~(in[919] ^ in[982]); 
    assign layer_0[8115] = ~in[150]; 
    assign layer_0[8116] = ~(in[610] | in[751]); 
    assign layer_0[8117] = in[106] & in[5]; 
    assign layer_0[8118] = ~in[494]; 
    assign layer_0[8119] = ~in[4] | (in[4] & in[644]); 
    assign layer_0[8120] = ~in[455] | (in[455] & in[744]); 
    assign layer_0[8121] = in[947] & ~in[997]; 
    assign layer_0[8122] = in[44] & in[724]; 
    assign layer_0[8123] = in[876] & ~in[984]; 
    assign layer_0[8124] = in[937] ^ in[699]; 
    assign layer_0[8125] = in[706] & ~in[430]; 
    assign layer_0[8126] = ~(in[618] ^ in[690]); 
    assign layer_0[8127] = ~in[619] | (in[619] & in[886]); 
    assign layer_0[8128] = in[97] & in[68]; 
    assign layer_0[8129] = in[78]; 
    assign layer_0[8130] = ~(in[774] & in[162]); 
    assign layer_0[8131] = ~in[924] | (in[895] & in[924]); 
    assign layer_0[8132] = in[232] ^ in[573]; 
    assign layer_0[8133] = in[213] ^ in[860]; 
    assign layer_0[8134] = in[318] | in[934]; 
    assign layer_0[8135] = in[724] & ~in[841]; 
    assign layer_0[8136] = in[417] ^ in[746]; 
    assign layer_0[8137] = in[570] & ~in[734]; 
    assign layer_0[8138] = ~(in[597] ^ in[161]); 
    assign layer_0[8139] = in[730] & ~in[740]; 
    assign layer_0[8140] = ~(in[765] | in[572]); 
    assign layer_0[8141] = in[953] & ~in[489]; 
    assign layer_0[8142] = ~(in[1000] | in[942]); 
    assign layer_0[8143] = in[461] & in[93]; 
    assign layer_0[8144] = in[937] | in[206]; 
    assign layer_0[8145] = ~(in[950] ^ in[596]); 
    assign layer_0[8146] = ~(in[61] | in[785]); 
    assign layer_0[8147] = in[549]; 
    assign layer_0[8148] = ~in[978] | (in[978] & in[240]); 
    assign layer_0[8149] = ~in[711]; 
    assign layer_0[8150] = ~in[718]; 
    assign layer_0[8151] = ~(in[603] ^ in[925]); 
    assign layer_0[8152] = ~(in[472] ^ in[245]); 
    assign layer_0[8153] = ~in[731]; 
    assign layer_0[8154] = ~(in[483] | in[34]); 
    assign layer_0[8155] = in[906] ^ in[943]; 
    assign layer_0[8156] = ~in[825]; 
    assign layer_0[8157] = in[1017] & ~in[273]; 
    assign layer_0[8158] = in[723] ^ in[435]; 
    assign layer_0[8159] = ~in[730] | (in[486] & in[730]); 
    assign layer_0[8160] = ~in[174]; 
    assign layer_0[8161] = in[607] ^ in[570]; 
    assign layer_0[8162] = ~(in[610] ^ in[674]); 
    assign layer_0[8163] = in[981] ^ in[675]; 
    assign layer_0[8164] = in[518] ^ in[519]; 
    assign layer_0[8165] = ~in[331] | (in[331] & in[95]); 
    assign layer_0[8166] = ~(in[149] ^ in[648]); 
    assign layer_0[8167] = in[1016]; 
    assign layer_0[8168] = in[1015] ^ in[789]; 
    assign layer_0[8169] = in[148]; 
    assign layer_0[8170] = ~(in[984] ^ in[774]); 
    assign layer_0[8171] = in[550] & in[550]; 
    assign layer_0[8172] = ~(in[664] ^ in[888]); 
    assign layer_0[8173] = in[653] ^ in[50]; 
    assign layer_0[8174] = ~in[552]; 
    assign layer_0[8175] = ~in[275] | (in[160] & in[275]); 
    assign layer_0[8176] = in[631] ^ in[632]; 
    assign layer_0[8177] = in[545] & ~in[342]; 
    assign layer_0[8178] = in[613] & ~in[242]; 
    assign layer_0[8179] = in[824]; 
    assign layer_0[8180] = ~(in[81] ^ in[533]); 
    assign layer_0[8181] = in[183] & in[488]; 
    assign layer_0[8182] = ~(in[787] & in[775]); 
    assign layer_0[8183] = ~(in[684] ^ in[564]); 
    assign layer_0[8184] = ~in[189] | (in[189] & in[565]); 
    assign layer_0[8185] = 1'b1; 
    assign layer_0[8186] = in[1005] ^ in[596]; 
    assign layer_0[8187] = in[206] ^ in[411]; 
    assign layer_0[8188] = ~in[866]; 
    assign layer_0[8189] = in[359] & ~in[952]; 
    assign layer_0[8190] = ~(in[239] | in[759]); 
    assign layer_0[8191] = 1'b0; 
    assign layer_0[8192] = in[12] & in[538]; 
    assign layer_0[8193] = ~in[632]; 
    assign layer_0[8194] = ~(in[10] ^ in[40]); 
    assign layer_0[8195] = in[963] | in[3]; 
    assign layer_0[8196] = ~in[629] | (in[757] & in[629]); 
    assign layer_0[8197] = in[209] ^ in[847]; 
    assign layer_0[8198] = in[367]; 
    assign layer_0[8199] = ~in[701] | (in[701] & in[790]); 
    assign layer_0[8200] = ~(in[651] | in[728]); 
    assign layer_0[8201] = ~(in[416] ^ in[476]); 
    assign layer_0[8202] = ~(in[776] | in[595]); 
    assign layer_0[8203] = ~(in[65] ^ in[539]); 
    assign layer_0[8204] = in[712] & ~in[976]; 
    assign layer_0[8205] = ~in[260] | (in[260] & in[679]); 
    assign layer_0[8206] = ~in[24] | (in[24] & in[284]); 
    assign layer_0[8207] = in[184] & in[189]; 
    assign layer_0[8208] = ~(in[323] ^ in[985]); 
    assign layer_0[8209] = in[8]; 
    assign layer_0[8210] = ~(in[367] ^ in[898]); 
    assign layer_0[8211] = ~in[789]; 
    assign layer_0[8212] = ~(in[18] | in[332]); 
    assign layer_0[8213] = in[485] ^ in[597]; 
    assign layer_0[8214] = in[596] ^ in[710]; 
    assign layer_0[8215] = in[177]; 
    assign layer_0[8216] = in[689] ^ in[76]; 
    assign layer_0[8217] = ~(in[35] ^ in[747]); 
    assign layer_0[8218] = ~(in[791] ^ in[696]); 
    assign layer_0[8219] = ~in[316]; 
    assign layer_0[8220] = ~(in[307] ^ in[792]); 
    assign layer_0[8221] = ~in[289]; 
    assign layer_0[8222] = ~in[243]; 
    assign layer_0[8223] = ~in[294] | (in[294] & in[533]); 
    assign layer_0[8224] = in[145] & ~in[449]; 
    assign layer_0[8225] = in[413]; 
    assign layer_0[8226] = ~(in[940] ^ in[563]); 
    assign layer_0[8227] = in[251] ^ in[500]; 
    assign layer_0[8228] = ~(in[59] ^ in[217]); 
    assign layer_0[8229] = in[536] & in[349]; 
    assign layer_0[8230] = 1'b1; 
    assign layer_0[8231] = ~in[378] | (in[627] & in[378]); 
    assign layer_0[8232] = in[428] & in[4]; 
    assign layer_0[8233] = in[858]; 
    assign layer_0[8234] = ~in[804]; 
    assign layer_0[8235] = ~in[944]; 
    assign layer_0[8236] = ~in[312]; 
    assign layer_0[8237] = in[643] ^ in[731]; 
    assign layer_0[8238] = in[962] ^ in[877]; 
    assign layer_0[8239] = ~(in[968] ^ in[21]); 
    assign layer_0[8240] = 1'b0; 
    assign layer_0[8241] = ~(in[503] & in[805]); 
    assign layer_0[8242] = in[110] ^ in[437]; 
    assign layer_0[8243] = ~in[888] | (in[754] & in[888]); 
    assign layer_0[8244] = in[704] ^ in[613]; 
    assign layer_0[8245] = ~(in[957] ^ in[703]); 
    assign layer_0[8246] = in[760]; 
    assign layer_0[8247] = in[806] ^ in[807]; 
    assign layer_0[8248] = in[29]; 
    assign layer_0[8249] = ~(in[644] | in[497]); 
    assign layer_0[8250] = ~(in[328] & in[398]); 
    assign layer_0[8251] = in[663]; 
    assign layer_0[8252] = in[341] & ~in[624]; 
    assign layer_0[8253] = ~in[80]; 
    assign layer_0[8254] = in[599] & ~in[311]; 
    assign layer_0[8255] = in[711]; 
    assign layer_0[8256] = ~in[956] | (in[996] & in[956]); 
    assign layer_0[8257] = ~(in[917] | in[190]); 
    assign layer_0[8258] = in[53]; 
    assign layer_0[8259] = ~(in[130] ^ in[301]); 
    assign layer_0[8260] = ~in[1]; 
    assign layer_0[8261] = ~in[985] | (in[985] & in[872]); 
    assign layer_0[8262] = ~(in[843] ^ in[667]); 
    assign layer_0[8263] = ~(in[695] ^ in[264]); 
    assign layer_0[8264] = ~(in[501] & in[781]); 
    assign layer_0[8265] = in[718] | in[874]; 
    assign layer_0[8266] = ~(in[571] ^ in[268]); 
    assign layer_0[8267] = in[396] | in[917]; 
    assign layer_0[8268] = in[261] ^ in[1011]; 
    assign layer_0[8269] = in[600] | in[45]; 
    assign layer_0[8270] = in[739] & in[728]; 
    assign layer_0[8271] = in[354]; 
    assign layer_0[8272] = in[759] ^ in[3]; 
    assign layer_0[8273] = in[539] ^ in[776]; 
    assign layer_0[8274] = ~in[362] | (in[362] & in[916]); 
    assign layer_0[8275] = in[517] & ~in[288]; 
    assign layer_0[8276] = in[198] ^ in[878]; 
    assign layer_0[8277] = ~(in[996] ^ in[629]); 
    assign layer_0[8278] = ~(in[970] & in[507]); 
    assign layer_0[8279] = 1'b0; 
    assign layer_0[8280] = ~in[821] | (in[821] & in[271]); 
    assign layer_0[8281] = ~in[920] | (in[920] & in[483]); 
    assign layer_0[8282] = ~in[578]; 
    assign layer_0[8283] = in[63] ^ in[607]; 
    assign layer_0[8284] = in[140]; 
    assign layer_0[8285] = in[235] ^ in[556]; 
    assign layer_0[8286] = ~in[538] | (in[951] & in[538]); 
    assign layer_0[8287] = ~in[776]; 
    assign layer_0[8288] = in[1016] ^ in[715]; 
    assign layer_0[8289] = in[212] & in[583]; 
    assign layer_0[8290] = in[320] & in[886]; 
    assign layer_0[8291] = in[252] & in[45]; 
    assign layer_0[8292] = ~in[503]; 
    assign layer_0[8293] = in[461]; 
    assign layer_0[8294] = in[194] & ~in[871]; 
    assign layer_0[8295] = ~(in[177] ^ in[397]); 
    assign layer_0[8296] = ~(in[856] | in[531]); 
    assign layer_0[8297] = ~in[859] | (in[859] & in[321]); 
    assign layer_0[8298] = in[551] & ~in[734]; 
    assign layer_0[8299] = ~in[299]; 
    assign layer_0[8300] = ~(in[917] ^ in[965]); 
    assign layer_0[8301] = ~(in[779] | in[729]); 
    assign layer_0[8302] = ~(in[612] ^ in[971]); 
    assign layer_0[8303] = in[491] & ~in[897]; 
    assign layer_0[8304] = ~(in[705] ^ in[583]); 
    assign layer_0[8305] = ~in[400]; 
    assign layer_0[8306] = in[838] & ~in[638]; 
    assign layer_0[8307] = in[703] ^ in[712]; 
    assign layer_0[8308] = in[645]; 
    assign layer_0[8309] = in[493] ^ in[844]; 
    assign layer_0[8310] = ~(in[275] ^ in[967]); 
    assign layer_0[8311] = in[837] | in[838]; 
    assign layer_0[8312] = ~(in[483] ^ in[716]); 
    assign layer_0[8313] = in[611] ^ in[807]; 
    assign layer_0[8314] = ~(in[884] ^ in[1007]); 
    assign layer_0[8315] = in[874] | in[346]; 
    assign layer_0[8316] = ~(in[628] ^ in[716]); 
    assign layer_0[8317] = in[689] & ~in[1003]; 
    assign layer_0[8318] = ~(in[627] ^ in[206]); 
    assign layer_0[8319] = in[283] ^ in[500]; 
    assign layer_0[8320] = ~(in[705] & in[85]); 
    assign layer_0[8321] = ~(in[551] ^ in[12]); 
    assign layer_0[8322] = in[984]; 
    assign layer_0[8323] = in[8] & ~in[517]; 
    assign layer_0[8324] = in[598]; 
    assign layer_0[8325] = ~in[904]; 
    assign layer_0[8326] = ~in[806]; 
    assign layer_0[8327] = ~in[263] | (in[522] & in[263]); 
    assign layer_0[8328] = ~(in[739] & in[741]); 
    assign layer_0[8329] = in[280] & in[500]; 
    assign layer_0[8330] = in[297] & ~in[343]; 
    assign layer_0[8331] = ~in[1002] | (in[1002] & in[33]); 
    assign layer_0[8332] = 1'b1; 
    assign layer_0[8333] = in[567]; 
    assign layer_0[8334] = ~(in[141] & in[242]); 
    assign layer_0[8335] = in[583] & ~in[801]; 
    assign layer_0[8336] = in[576]; 
    assign layer_0[8337] = ~in[261]; 
    assign layer_0[8338] = in[365] | in[904]; 
    assign layer_0[8339] = ~in[867]; 
    assign layer_0[8340] = in[266] | in[448]; 
    assign layer_0[8341] = ~(in[831] & in[527]); 
    assign layer_0[8342] = in[650] & in[366]; 
    assign layer_0[8343] = ~(in[971] & in[442]); 
    assign layer_0[8344] = in[490] & in[147]; 
    assign layer_0[8345] = ~in[307]; 
    assign layer_0[8346] = ~(in[546] | in[372]); 
    assign layer_0[8347] = in[615] & ~in[552]; 
    assign layer_0[8348] = ~in[252]; 
    assign layer_0[8349] = in[97] & ~in[885]; 
    assign layer_0[8350] = ~(in[677] ^ in[356]); 
    assign layer_0[8351] = in[140] & ~in[412]; 
    assign layer_0[8352] = in[699] ^ in[611]; 
    assign layer_0[8353] = in[372] & in[283]; 
    assign layer_0[8354] = in[752] | in[951]; 
    assign layer_0[8355] = in[657] ^ in[22]; 
    assign layer_0[8356] = ~(in[340] | in[713]); 
    assign layer_0[8357] = in[795] | in[65]; 
    assign layer_0[8358] = ~(in[764] ^ in[308]); 
    assign layer_0[8359] = in[690] & ~in[912]; 
    assign layer_0[8360] = in[936] ^ in[401]; 
    assign layer_0[8361] = in[911]; 
    assign layer_0[8362] = ~(in[597] ^ in[62]); 
    assign layer_0[8363] = ~(in[129] & in[23]); 
    assign layer_0[8364] = in[333] ^ in[429]; 
    assign layer_0[8365] = ~(in[924] | in[700]); 
    assign layer_0[8366] = ~in[549]; 
    assign layer_0[8367] = in[265] ^ in[402]; 
    assign layer_0[8368] = ~(in[619] ^ in[98]); 
    assign layer_0[8369] = in[239] ^ in[6]; 
    assign layer_0[8370] = in[46]; 
    assign layer_0[8371] = ~(in[1014] | in[109]); 
    assign layer_0[8372] = ~(in[596] & in[791]); 
    assign layer_0[8373] = in[69] | in[977]; 
    assign layer_0[8374] = ~(in[76] | in[458]); 
    assign layer_0[8375] = in[747] ^ in[516]; 
    assign layer_0[8376] = in[319] & ~in[985]; 
    assign layer_0[8377] = ~in[597] | (in[597] & in[997]); 
    assign layer_0[8378] = ~in[113] | (in[305] & in[113]); 
    assign layer_0[8379] = ~(in[714] ^ in[957]); 
    assign layer_0[8380] = in[888] ^ in[889]; 
    assign layer_0[8381] = in[623] ^ in[327]; 
    assign layer_0[8382] = in[308] ^ in[258]; 
    assign layer_0[8383] = in[493] ^ in[892]; 
    assign layer_0[8384] = ~(in[464] ^ in[296]); 
    assign layer_0[8385] = in[245] ^ in[522]; 
    assign layer_0[8386] = in[7] | in[31]; 
    assign layer_0[8387] = in[933] & ~in[776]; 
    assign layer_0[8388] = ~(in[942] ^ in[241]); 
    assign layer_0[8389] = ~(in[554] ^ in[388]); 
    assign layer_0[8390] = in[811] & in[342]; 
    assign layer_0[8391] = in[555] ^ in[886]; 
    assign layer_0[8392] = ~in[263] | (in[505] & in[263]); 
    assign layer_0[8393] = in[94]; 
    assign layer_0[8394] = ~(in[100] | in[544]); 
    assign layer_0[8395] = ~(in[846] ^ in[700]); 
    assign layer_0[8396] = in[361] & in[860]; 
    assign layer_0[8397] = in[552] | in[98]; 
    assign layer_0[8398] = in[839] ^ in[971]; 
    assign layer_0[8399] = ~in[709] | (in[584] & in[709]); 
    assign layer_0[8400] = in[827] ^ in[286]; 
    assign layer_0[8401] = ~in[36] | (in[36] & in[607]); 
    assign layer_0[8402] = in[291] ^ in[263]; 
    assign layer_0[8403] = in[279] ^ in[840]; 
    assign layer_0[8404] = in[697] & in[614]; 
    assign layer_0[8405] = in[75] ^ in[795]; 
    assign layer_0[8406] = ~(in[951] ^ in[952]); 
    assign layer_0[8407] = ~(in[998] ^ in[999]); 
    assign layer_0[8408] = ~in[240]; 
    assign layer_0[8409] = in[775] ^ in[748]; 
    assign layer_0[8410] = ~(in[660] ^ in[741]); 
    assign layer_0[8411] = in[429] & ~in[944]; 
    assign layer_0[8412] = ~(in[92] ^ in[636]); 
    assign layer_0[8413] = ~(in[266] ^ in[910]); 
    assign layer_0[8414] = ~in[532]; 
    assign layer_0[8415] = in[993] ^ in[590]; 
    assign layer_0[8416] = in[466] ^ in[129]; 
    assign layer_0[8417] = ~(in[900] ^ in[1006]); 
    assign layer_0[8418] = ~(in[698] ^ in[700]); 
    assign layer_0[8419] = ~(in[698] ^ in[826]); 
    assign layer_0[8420] = in[811] | in[859]; 
    assign layer_0[8421] = in[728] & ~in[747]; 
    assign layer_0[8422] = ~(in[904] ^ in[252]); 
    assign layer_0[8423] = ~in[262] | (in[468] & in[262]); 
    assign layer_0[8424] = in[181] | in[867]; 
    assign layer_0[8425] = in[868] ^ in[453]; 
    assign layer_0[8426] = in[748] ^ in[956]; 
    assign layer_0[8427] = ~(in[259] ^ in[746]); 
    assign layer_0[8428] = in[160] & ~in[98]; 
    assign layer_0[8429] = ~(in[260] ^ in[870]); 
    assign layer_0[8430] = ~(in[618] & in[325]); 
    assign layer_0[8431] = ~in[95]; 
    assign layer_0[8432] = ~in[465] | (in[692] & in[465]); 
    assign layer_0[8433] = in[357] & ~in[302]; 
    assign layer_0[8434] = ~in[371]; 
    assign layer_0[8435] = in[111] ^ in[731]; 
    assign layer_0[8436] = ~(in[843] ^ in[2]); 
    assign layer_0[8437] = ~in[390] | (in[504] & in[390]); 
    assign layer_0[8438] = in[126] & in[39]; 
    assign layer_0[8439] = in[872] ^ in[955]; 
    assign layer_0[8440] = ~in[80]; 
    assign layer_0[8441] = ~in[292]; 
    assign layer_0[8442] = ~in[663] | (in[663] & in[21]); 
    assign layer_0[8443] = ~in[1002] | (in[1002] & in[838]); 
    assign layer_0[8444] = ~(in[856] ^ in[898]); 
    assign layer_0[8445] = ~in[872]; 
    assign layer_0[8446] = in[759]; 
    assign layer_0[8447] = ~(in[450] ^ in[342]); 
    assign layer_0[8448] = ~in[409] | (in[980] & in[409]); 
    assign layer_0[8449] = in[640] ^ in[473]; 
    assign layer_0[8450] = in[487] ^ in[569]; 
    assign layer_0[8451] = ~(in[572] | in[873]); 
    assign layer_0[8452] = ~(in[867] & in[556]); 
    assign layer_0[8453] = in[94]; 
    assign layer_0[8454] = ~(in[517] | in[540]); 
    assign layer_0[8455] = in[684] ^ in[113]; 
    assign layer_0[8456] = ~(in[350] ^ in[463]); 
    assign layer_0[8457] = in[101] | in[783]; 
    assign layer_0[8458] = ~(in[603] & in[135]); 
    assign layer_0[8459] = in[921] ^ in[381]; 
    assign layer_0[8460] = ~in[954]; 
    assign layer_0[8461] = ~(in[161] | in[371]); 
    assign layer_0[8462] = ~(in[150] & in[823]); 
    assign layer_0[8463] = in[264] ^ in[487]; 
    assign layer_0[8464] = in[930] | in[555]; 
    assign layer_0[8465] = ~(in[1018] & in[376]); 
    assign layer_0[8466] = in[548] ^ in[900]; 
    assign layer_0[8467] = in[778] | in[798]; 
    assign layer_0[8468] = in[66]; 
    assign layer_0[8469] = in[428] ^ in[371]; 
    assign layer_0[8470] = in[19] ^ in[78]; 
    assign layer_0[8471] = in[699]; 
    assign layer_0[8472] = ~(in[277] | in[176]); 
    assign layer_0[8473] = ~(in[627] & in[450]); 
    assign layer_0[8474] = in[356] ^ in[249]; 
    assign layer_0[8475] = ~in[492]; 
    assign layer_0[8476] = in[253] ^ in[902]; 
    assign layer_0[8477] = in[623] ^ in[494]; 
    assign layer_0[8478] = ~(in[808] ^ in[806]); 
    assign layer_0[8479] = in[839] ^ in[184]; 
    assign layer_0[8480] = ~in[587]; 
    assign layer_0[8481] = in[778] ^ in[243]; 
    assign layer_0[8482] = ~in[241]; 
    assign layer_0[8483] = in[522] & ~in[916]; 
    assign layer_0[8484] = in[714] ^ in[968]; 
    assign layer_0[8485] = in[960]; 
    assign layer_0[8486] = ~(in[18] ^ in[516]); 
    assign layer_0[8487] = in[871] ^ in[926]; 
    assign layer_0[8488] = 1'b1; 
    assign layer_0[8489] = in[854] ^ in[692]; 
    assign layer_0[8490] = ~in[603] | (in[859] & in[603]); 
    assign layer_0[8491] = ~in[292]; 
    assign layer_0[8492] = ~(in[886] ^ in[901]); 
    assign layer_0[8493] = in[350]; 
    assign layer_0[8494] = 1'b1; 
    assign layer_0[8495] = in[807] & in[522]; 
    assign layer_0[8496] = ~in[244] | (in[244] & in[107]); 
    assign layer_0[8497] = in[279] & ~in[756]; 
    assign layer_0[8498] = ~in[592] | (in[91] & in[592]); 
    assign layer_0[8499] = ~in[898] | (in[898] & in[596]); 
    assign layer_0[8500] = in[114] & in[53]; 
    assign layer_0[8501] = in[874]; 
    assign layer_0[8502] = ~(in[270] | in[1016]); 
    assign layer_0[8503] = in[583] & ~in[297]; 
    assign layer_0[8504] = ~(in[614] | in[738]); 
    assign layer_0[8505] = in[723] & ~in[551]; 
    assign layer_0[8506] = ~(in[807] ^ in[242]); 
    assign layer_0[8507] = in[372] & ~in[640]; 
    assign layer_0[8508] = ~(in[546] & in[787]); 
    assign layer_0[8509] = in[699] ^ in[885]; 
    assign layer_0[8510] = ~(in[807] ^ in[1000]); 
    assign layer_0[8511] = ~(in[403] ^ in[869]); 
    assign layer_0[8512] = in[476] ^ in[213]; 
    assign layer_0[8513] = ~(in[537] | in[285]); 
    assign layer_0[8514] = ~(in[751] & in[352]); 
    assign layer_0[8515] = in[321]; 
    assign layer_0[8516] = in[921] ^ in[533]; 
    assign layer_0[8517] = in[28] & ~in[333]; 
    assign layer_0[8518] = in[708] ^ in[466]; 
    assign layer_0[8519] = ~(in[129] & in[460]); 
    assign layer_0[8520] = ~(in[191] | in[1010]); 
    assign layer_0[8521] = ~(in[70] ^ in[224]); 
    assign layer_0[8522] = in[3] & in[989]; 
    assign layer_0[8523] = in[907] ^ in[562]; 
    assign layer_0[8524] = in[715] & ~in[885]; 
    assign layer_0[8525] = in[581] & ~in[685]; 
    assign layer_0[8526] = ~(in[871] & in[957]); 
    assign layer_0[8527] = ~(in[370] ^ in[538]); 
    assign layer_0[8528] = ~(in[549] ^ in[370]); 
    assign layer_0[8529] = ~in[371] | (in[965] & in[371]); 
    assign layer_0[8530] = ~in[401] | (in[401] & in[564]); 
    assign layer_0[8531] = in[134] & in[375]; 
    assign layer_0[8532] = in[871] ^ in[888]; 
    assign layer_0[8533] = ~(in[64] & in[309]); 
    assign layer_0[8534] = ~in[585] | (in[764] & in[585]); 
    assign layer_0[8535] = in[533] ^ in[981]; 
    assign layer_0[8536] = in[497] | in[879]; 
    assign layer_0[8537] = in[7] & ~in[519]; 
    assign layer_0[8538] = in[454] ^ in[907]; 
    assign layer_0[8539] = ~(in[761] ^ in[793]); 
    assign layer_0[8540] = ~(in[885] | in[901]); 
    assign layer_0[8541] = ~(in[583] ^ in[870]); 
    assign layer_0[8542] = ~(in[426] ^ in[267]); 
    assign layer_0[8543] = in[889] & ~in[854]; 
    assign layer_0[8544] = in[698]; 
    assign layer_0[8545] = ~in[553] | (in[210] & in[553]); 
    assign layer_0[8546] = ~(in[746] ^ in[337]); 
    assign layer_0[8547] = in[936] & ~in[854]; 
    assign layer_0[8548] = ~in[735] | (in[735] & in[773]); 
    assign layer_0[8549] = in[957] & ~in[573]; 
    assign layer_0[8550] = ~(in[267] ^ in[271]); 
    assign layer_0[8551] = ~(in[728] ^ in[157]); 
    assign layer_0[8552] = in[859] ^ in[790]; 
    assign layer_0[8553] = in[734] | in[797]; 
    assign layer_0[8554] = in[922] ^ in[508]; 
    assign layer_0[8555] = in[366] & ~in[739]; 
    assign layer_0[8556] = in[705]; 
    assign layer_0[8557] = in[823] ^ in[449]; 
    assign layer_0[8558] = in[301] | in[793]; 
    assign layer_0[8559] = in[355]; 
    assign layer_0[8560] = ~(in[601] & in[475]); 
    assign layer_0[8561] = in[95] & ~in[840]; 
    assign layer_0[8562] = ~in[999]; 
    assign layer_0[8563] = ~(in[839] ^ in[990]); 
    assign layer_0[8564] = ~(in[500] ^ in[1015]); 
    assign layer_0[8565] = in[460] & ~in[525]; 
    assign layer_0[8566] = in[487]; 
    assign layer_0[8567] = in[892] & in[634]; 
    assign layer_0[8568] = ~(in[340] & in[396]); 
    assign layer_0[8569] = in[449] & ~in[981]; 
    assign layer_0[8570] = ~(in[351] ^ in[453]); 
    assign layer_0[8571] = ~(in[365] & in[746]); 
    assign layer_0[8572] = ~(in[748] ^ in[261]); 
    assign layer_0[8573] = ~in[822] | (in[822] & in[948]); 
    assign layer_0[8574] = ~(in[52] ^ in[20]); 
    assign layer_0[8575] = in[522] ^ in[614]; 
    assign layer_0[8576] = ~in[538] | (in[7] & in[538]); 
    assign layer_0[8577] = ~(in[563] ^ in[473]); 
    assign layer_0[8578] = in[565] & ~in[279]; 
    assign layer_0[8579] = in[616] & in[296]; 
    assign layer_0[8580] = ~in[971] | (in[971] & in[796]); 
    assign layer_0[8581] = ~in[623] | (in[578] & in[623]); 
    assign layer_0[8582] = ~(in[445] & in[296]); 
    assign layer_0[8583] = ~(in[953] ^ in[952]); 
    assign layer_0[8584] = ~(in[827] | in[790]); 
    assign layer_0[8585] = ~(in[992] | in[944]); 
    assign layer_0[8586] = in[810] | in[793]; 
    assign layer_0[8587] = in[612] ^ in[251]; 
    assign layer_0[8588] = in[57]; 
    assign layer_0[8589] = in[878]; 
    assign layer_0[8590] = in[147]; 
    assign layer_0[8591] = in[984] ^ in[982]; 
    assign layer_0[8592] = ~(in[968] & in[709]); 
    assign layer_0[8593] = in[818]; 
    assign layer_0[8594] = ~in[727]; 
    assign layer_0[8595] = ~in[565] | (in[890] & in[565]); 
    assign layer_0[8596] = in[210] ^ in[98]; 
    assign layer_0[8597] = ~(in[158] & in[989]); 
    assign layer_0[8598] = in[253] & ~in[418]; 
    assign layer_0[8599] = ~in[909] | (in[909] & in[557]); 
    assign layer_0[8600] = in[156] & in[654]; 
    assign layer_0[8601] = in[693] ^ in[366]; 
    assign layer_0[8602] = in[845] & ~in[930]; 
    assign layer_0[8603] = in[691] | in[466]; 
    assign layer_0[8604] = in[996]; 
    assign layer_0[8605] = in[193] ^ in[111]; 
    assign layer_0[8606] = ~(in[523] & in[218]); 
    assign layer_0[8607] = ~(in[537] & in[534]); 
    assign layer_0[8608] = ~(in[382] ^ in[521]); 
    assign layer_0[8609] = in[647] ^ in[890]; 
    assign layer_0[8610] = in[612] & in[332]; 
    assign layer_0[8611] = ~(in[414] ^ in[700]); 
    assign layer_0[8612] = 1'b0; 
    assign layer_0[8613] = in[251] & ~in[788]; 
    assign layer_0[8614] = in[825]; 
    assign layer_0[8615] = in[533] ^ in[519]; 
    assign layer_0[8616] = 1'b1; 
    assign layer_0[8617] = ~in[845] | (in[845] & in[966]); 
    assign layer_0[8618] = ~(in[33] | in[518]); 
    assign layer_0[8619] = in[632] & in[427]; 
    assign layer_0[8620] = in[870] & in[621]; 
    assign layer_0[8621] = in[54] ^ in[651]; 
    assign layer_0[8622] = ~in[925] | (in[925] & in[735]); 
    assign layer_0[8623] = ~(in[67] & in[491]); 
    assign layer_0[8624] = in[844] ^ in[1005]; 
    assign layer_0[8625] = ~(in[921] ^ in[218]); 
    assign layer_0[8626] = ~(in[123] ^ in[642]); 
    assign layer_0[8627] = in[835] & in[365]; 
    assign layer_0[8628] = in[264] & ~in[763]; 
    assign layer_0[8629] = ~in[595]; 
    assign layer_0[8630] = in[664] ^ in[989]; 
    assign layer_0[8631] = in[446] ^ in[334]; 
    assign layer_0[8632] = ~(in[947] ^ in[795]); 
    assign layer_0[8633] = in[260] & ~in[598]; 
    assign layer_0[8634] = in[189]; 
    assign layer_0[8635] = in[227] & ~in[733]; 
    assign layer_0[8636] = ~(in[13] ^ in[21]); 
    assign layer_0[8637] = ~(in[195] & in[775]); 
    assign layer_0[8638] = in[264] & ~in[789]; 
    assign layer_0[8639] = ~(in[432] ^ in[489]); 
    assign layer_0[8640] = ~(in[1018] ^ in[366]); 
    assign layer_0[8641] = in[604] ^ in[254]; 
    assign layer_0[8642] = in[639] ^ in[950]; 
    assign layer_0[8643] = ~(in[61] ^ in[950]); 
    assign layer_0[8644] = ~in[598] | (in[160] & in[598]); 
    assign layer_0[8645] = in[873] ^ in[520]; 
    assign layer_0[8646] = in[26]; 
    assign layer_0[8647] = ~in[387]; 
    assign layer_0[8648] = in[568]; 
    assign layer_0[8649] = in[995]; 
    assign layer_0[8650] = in[144] & in[394]; 
    assign layer_0[8651] = ~in[90] | (in[90] & in[941]); 
    assign layer_0[8652] = ~in[497] | (in[905] & in[497]); 
    assign layer_0[8653] = ~in[746] | (in[746] & in[503]); 
    assign layer_0[8654] = in[618] ^ in[599]; 
    assign layer_0[8655] = ~(in[445] & in[38]); 
    assign layer_0[8656] = in[678] ^ in[264]; 
    assign layer_0[8657] = in[588] ^ in[477]; 
    assign layer_0[8658] = ~in[256]; 
    assign layer_0[8659] = ~(in[890] ^ in[648]); 
    assign layer_0[8660] = ~(in[487] ^ in[141]); 
    assign layer_0[8661] = in[299] ^ in[985]; 
    assign layer_0[8662] = in[37] & ~in[570]; 
    assign layer_0[8663] = ~in[708]; 
    assign layer_0[8664] = ~(in[592] | in[771]); 
    assign layer_0[8665] = in[712] & ~in[902]; 
    assign layer_0[8666] = ~in[193] | (in[766] & in[193]); 
    assign layer_0[8667] = in[342] ^ in[356]; 
    assign layer_0[8668] = in[569]; 
    assign layer_0[8669] = in[806] ^ in[971]; 
    assign layer_0[8670] = in[433] | in[240]; 
    assign layer_0[8671] = in[682] & ~in[790]; 
    assign layer_0[8672] = ~(in[826] ^ in[569]); 
    assign layer_0[8673] = ~(in[631] | in[498]); 
    assign layer_0[8674] = ~in[184] | (in[184] & in[835]); 
    assign layer_0[8675] = ~in[875] | (in[875] & in[573]); 
    assign layer_0[8676] = in[889] & in[979]; 
    assign layer_0[8677] = in[984] | in[888]; 
    assign layer_0[8678] = in[98] ^ in[555]; 
    assign layer_0[8679] = ~(in[318] | in[4]); 
    assign layer_0[8680] = ~(in[744] ^ in[715]); 
    assign layer_0[8681] = ~(in[669] & in[838]); 
    assign layer_0[8682] = in[714]; 
    assign layer_0[8683] = in[611] ^ in[485]; 
    assign layer_0[8684] = ~in[275]; 
    assign layer_0[8685] = ~in[131] | (in[131] & in[999]); 
    assign layer_0[8686] = in[681] & ~in[997]; 
    assign layer_0[8687] = in[661] ^ in[981]; 
    assign layer_0[8688] = ~in[20] | (in[20] & in[268]); 
    assign layer_0[8689] = ~in[252] | (in[252] & in[763]); 
    assign layer_0[8690] = ~(in[663] & in[666]); 
    assign layer_0[8691] = ~(in[176] | in[935]); 
    assign layer_0[8692] = ~(in[476] ^ in[667]); 
    assign layer_0[8693] = ~in[179] | (in[179] & in[809]); 
    assign layer_0[8694] = ~(in[630] ^ in[934]); 
    assign layer_0[8695] = ~(in[33] ^ in[503]); 
    assign layer_0[8696] = ~(in[444] ^ in[333]); 
    assign layer_0[8697] = ~(in[306] ^ in[163]); 
    assign layer_0[8698] = in[594] | in[422]; 
    assign layer_0[8699] = ~(in[454] & in[912]); 
    assign layer_0[8700] = ~in[297] | (in[297] & in[321]); 
    assign layer_0[8701] = ~in[934]; 
    assign layer_0[8702] = in[697] & in[136]; 
    assign layer_0[8703] = ~in[40]; 
    assign layer_0[8704] = ~(in[413] ^ in[356]); 
    assign layer_0[8705] = in[273] | in[597]; 
    assign layer_0[8706] = in[580]; 
    assign layer_0[8707] = ~(in[552] ^ in[467]); 
    assign layer_0[8708] = ~in[884]; 
    assign layer_0[8709] = in[521] & ~in[365]; 
    assign layer_0[8710] = ~in[1002] | (in[1002] & in[790]); 
    assign layer_0[8711] = in[931] & in[430]; 
    assign layer_0[8712] = in[981] | in[847]; 
    assign layer_0[8713] = in[624] | in[669]; 
    assign layer_0[8714] = ~(in[889] ^ in[953]); 
    assign layer_0[8715] = in[889] | in[1016]; 
    assign layer_0[8716] = in[946] ^ in[449]; 
    assign layer_0[8717] = in[821] & ~in[514]; 
    assign layer_0[8718] = ~(in[300] & in[243]); 
    assign layer_0[8719] = ~in[487]; 
    assign layer_0[8720] = ~(in[181] ^ in[589]); 
    assign layer_0[8721] = in[1015] | in[948]; 
    assign layer_0[8722] = in[518] | in[29]; 
    assign layer_0[8723] = ~(in[38] & in[179]); 
    assign layer_0[8724] = in[284]; 
    assign layer_0[8725] = in[347] & ~in[28]; 
    assign layer_0[8726] = in[808] ^ in[565]; 
    assign layer_0[8727] = ~(in[827] | in[807]); 
    assign layer_0[8728] = ~in[285]; 
    assign layer_0[8729] = ~in[886] | (in[756] & in[886]); 
    assign layer_0[8730] = ~in[993]; 
    assign layer_0[8731] = ~(in[505] & in[687]); 
    assign layer_0[8732] = in[925] ^ in[590]; 
    assign layer_0[8733] = in[651] & ~in[89]; 
    assign layer_0[8734] = in[39] & in[55]; 
    assign layer_0[8735] = in[675] & in[18]; 
    assign layer_0[8736] = ~in[252]; 
    assign layer_0[8737] = in[851]; 
    assign layer_0[8738] = in[323] | in[915]; 
    assign layer_0[8739] = ~(in[457] | in[910]); 
    assign layer_0[8740] = ~in[155] | (in[979] & in[155]); 
    assign layer_0[8741] = ~in[663]; 
    assign layer_0[8742] = in[948] | in[844]; 
    assign layer_0[8743] = ~in[214] | (in[825] & in[214]); 
    assign layer_0[8744] = ~in[139]; 
    assign layer_0[8745] = in[221] | in[715]; 
    assign layer_0[8746] = ~(in[874] | in[844]); 
    assign layer_0[8747] = ~(in[290] | in[612]); 
    assign layer_0[8748] = in[273] & in[682]; 
    assign layer_0[8749] = in[219] & ~in[12]; 
    assign layer_0[8750] = ~in[635] | (in[635] & in[1000]); 
    assign layer_0[8751] = ~in[153] | (in[595] & in[153]); 
    assign layer_0[8752] = in[969] & ~in[48]; 
    assign layer_0[8753] = ~(in[251] ^ in[479]); 
    assign layer_0[8754] = ~(in[206] ^ in[854]); 
    assign layer_0[8755] = in[341] & ~in[413]; 
    assign layer_0[8756] = ~in[360] | (in[360] & in[831]); 
    assign layer_0[8757] = in[537] ^ in[885]; 
    assign layer_0[8758] = in[394] ^ in[621]; 
    assign layer_0[8759] = in[613] ^ in[189]; 
    assign layer_0[8760] = in[587] ^ in[820]; 
    assign layer_0[8761] = ~in[28]; 
    assign layer_0[8762] = ~(in[533] & in[562]); 
    assign layer_0[8763] = ~in[485] | (in[485] & in[439]); 
    assign layer_0[8764] = in[788] | in[693]; 
    assign layer_0[8765] = in[299] & ~in[760]; 
    assign layer_0[8766] = in[477] & ~in[473]; 
    assign layer_0[8767] = in[182] & in[685]; 
    assign layer_0[8768] = in[262] ^ in[242]; 
    assign layer_0[8769] = in[846]; 
    assign layer_0[8770] = ~(in[569] ^ in[34]); 
    assign layer_0[8771] = in[806] & in[699]; 
    assign layer_0[8772] = ~in[297]; 
    assign layer_0[8773] = in[775] | in[541]; 
    assign layer_0[8774] = ~(in[492] & in[162]); 
    assign layer_0[8775] = ~in[49]; 
    assign layer_0[8776] = in[844] | in[524]; 
    assign layer_0[8777] = ~in[914]; 
    assign layer_0[8778] = in[930] ^ in[384]; 
    assign layer_0[8779] = ~in[841]; 
    assign layer_0[8780] = in[793] ^ in[792]; 
    assign layer_0[8781] = in[956] & in[730]; 
    assign layer_0[8782] = ~(in[365] ^ in[1003]); 
    assign layer_0[8783] = in[699]; 
    assign layer_0[8784] = ~in[81] | (in[961] & in[81]); 
    assign layer_0[8785] = ~(in[116] | in[525]); 
    assign layer_0[8786] = in[115] & ~in[1019]; 
    assign layer_0[8787] = ~(in[466] ^ in[856]); 
    assign layer_0[8788] = in[100] ^ in[648]; 
    assign layer_0[8789] = ~(in[901] ^ in[690]); 
    assign layer_0[8790] = in[786] & ~in[309]; 
    assign layer_0[8791] = in[600] ^ in[265]; 
    assign layer_0[8792] = in[522]; 
    assign layer_0[8793] = ~(in[647] ^ in[906]); 
    assign layer_0[8794] = in[838] & in[235]; 
    assign layer_0[8795] = in[740] & ~in[845]; 
    assign layer_0[8796] = in[523]; 
    assign layer_0[8797] = ~(in[129] | in[851]); 
    assign layer_0[8798] = in[217] | in[919]; 
    assign layer_0[8799] = in[669] ^ in[729]; 
    assign layer_0[8800] = in[763] | in[594]; 
    assign layer_0[8801] = in[1002] & ~in[194]; 
    assign layer_0[8802] = ~in[247]; 
    assign layer_0[8803] = ~(in[553] | in[839]); 
    assign layer_0[8804] = ~in[679]; 
    assign layer_0[8805] = ~(in[663] & in[87]); 
    assign layer_0[8806] = ~in[72] | (in[72] & in[749]); 
    assign layer_0[8807] = in[333] & ~in[742]; 
    assign layer_0[8808] = 1'b0; 
    assign layer_0[8809] = in[131] | in[999]; 
    assign layer_0[8810] = in[365] ^ in[476]; 
    assign layer_0[8811] = ~(in[947] ^ in[574]); 
    assign layer_0[8812] = in[99] | in[1014]; 
    assign layer_0[8813] = ~(in[454] & in[98]); 
    assign layer_0[8814] = ~(in[573] ^ in[44]); 
    assign layer_0[8815] = ~(in[973] | in[129]); 
    assign layer_0[8816] = ~(in[97] | in[723]); 
    assign layer_0[8817] = ~(in[950] ^ in[128]); 
    assign layer_0[8818] = ~(in[62] | in[270]); 
    assign layer_0[8819] = ~(in[185] | in[624]); 
    assign layer_0[8820] = ~(in[757] ^ in[669]); 
    assign layer_0[8821] = ~(in[538] | in[78]); 
    assign layer_0[8822] = in[489]; 
    assign layer_0[8823] = in[391] & in[311]; 
    assign layer_0[8824] = in[77] ^ in[660]; 
    assign layer_0[8825] = in[15]; 
    assign layer_0[8826] = in[465] ^ in[956]; 
    assign layer_0[8827] = ~in[20] | (in[20] & in[177]); 
    assign layer_0[8828] = ~(in[816] | in[872]); 
    assign layer_0[8829] = in[572] | in[661]; 
    assign layer_0[8830] = in[994] | in[633]; 
    assign layer_0[8831] = ~(in[179] ^ in[587]); 
    assign layer_0[8832] = in[841] ^ in[838]; 
    assign layer_0[8833] = ~(in[678] ^ in[939]); 
    assign layer_0[8834] = ~(in[587] ^ in[1015]); 
    assign layer_0[8835] = ~(in[290] ^ in[347]); 
    assign layer_0[8836] = in[823]; 
    assign layer_0[8837] = in[635] ^ in[5]; 
    assign layer_0[8838] = in[626] ^ in[206]; 
    assign layer_0[8839] = in[953] ^ in[951]; 
    assign layer_0[8840] = in[520] ^ in[387]; 
    assign layer_0[8841] = ~in[295]; 
    assign layer_0[8842] = ~(in[831] | in[373]); 
    assign layer_0[8843] = in[658] ^ in[537]; 
    assign layer_0[8844] = in[136] & in[134]; 
    assign layer_0[8845] = in[906] ^ in[591]; 
    assign layer_0[8846] = in[253] & ~in[111]; 
    assign layer_0[8847] = ~(in[910] ^ in[316]); 
    assign layer_0[8848] = in[792] ^ in[825]; 
    assign layer_0[8849] = in[942] ^ in[607]; 
    assign layer_0[8850] = ~in[262] | (in[556] & in[262]); 
    assign layer_0[8851] = ~(in[364] ^ in[918]); 
    assign layer_0[8852] = ~(in[888] ^ in[738]); 
    assign layer_0[8853] = ~in[575]; 
    assign layer_0[8854] = in[66]; 
    assign layer_0[8855] = in[464] ^ in[172]; 
    assign layer_0[8856] = 1'b0; 
    assign layer_0[8857] = ~in[1014] | (in[924] & in[1014]); 
    assign layer_0[8858] = in[176] | in[564]; 
    assign layer_0[8859] = in[853] ^ in[886]; 
    assign layer_0[8860] = in[854] & in[756]; 
    assign layer_0[8861] = ~in[568]; 
    assign layer_0[8862] = ~(in[855] | in[860]); 
    assign layer_0[8863] = in[977] ^ in[416]; 
    assign layer_0[8864] = in[683] & ~in[858]; 
    assign layer_0[8865] = ~(in[306] ^ in[202]); 
    assign layer_0[8866] = ~(in[606] ^ in[901]); 
    assign layer_0[8867] = in[23]; 
    assign layer_0[8868] = ~in[275]; 
    assign layer_0[8869] = ~in[875] | (in[875] & in[880]); 
    assign layer_0[8870] = in[692]; 
    assign layer_0[8871] = ~(in[7] & in[572]); 
    assign layer_0[8872] = ~in[534] | (in[534] & in[1004]); 
    assign layer_0[8873] = in[938] | in[768]; 
    assign layer_0[8874] = ~(in[553] ^ in[691]); 
    assign layer_0[8875] = in[905] | in[45]; 
    assign layer_0[8876] = in[355] & ~in[352]; 
    assign layer_0[8877] = in[701]; 
    assign layer_0[8878] = ~in[108] | (in[108] & in[471]); 
    assign layer_0[8879] = ~(in[885] & in[144]); 
    assign layer_0[8880] = ~in[13]; 
    assign layer_0[8881] = ~in[65] | (in[965] & in[65]); 
    assign layer_0[8882] = in[533]; 
    assign layer_0[8883] = in[233] & in[494]; 
    assign layer_0[8884] = ~(in[984] | in[163]); 
    assign layer_0[8885] = ~in[373]; 
    assign layer_0[8886] = ~(in[749] ^ in[929]); 
    assign layer_0[8887] = in[461] ^ in[260]; 
    assign layer_0[8888] = ~(in[449] ^ in[113]); 
    assign layer_0[8889] = in[541] & in[708]; 
    assign layer_0[8890] = ~(in[562] ^ in[550]); 
    assign layer_0[8891] = ~in[324] | (in[686] & in[324]); 
    assign layer_0[8892] = in[886] | in[5]; 
    assign layer_0[8893] = ~in[263]; 
    assign layer_0[8894] = in[907] & ~in[70]; 
    assign layer_0[8895] = in[664] & ~in[994]; 
    assign layer_0[8896] = ~(in[202] & in[477]); 
    assign layer_0[8897] = in[106] ^ in[754]; 
    assign layer_0[8898] = in[808]; 
    assign layer_0[8899] = ~(in[70] | in[827]); 
    assign layer_0[8900] = in[293]; 
    assign layer_0[8901] = in[860] ^ in[878]; 
    assign layer_0[8902] = in[537] | in[705]; 
    assign layer_0[8903] = ~in[672] | (in[607] & in[672]); 
    assign layer_0[8904] = ~in[196] | (in[196] & in[793]); 
    assign layer_0[8905] = ~(in[742] & in[19]); 
    assign layer_0[8906] = ~in[186] | (in[186] & in[310]); 
    assign layer_0[8907] = in[283] ^ in[906]; 
    assign layer_0[8908] = in[313] & in[936]; 
    assign layer_0[8909] = in[654]; 
    assign layer_0[8910] = in[836] | in[821]; 
    assign layer_0[8911] = ~in[378] | (in[943] & in[378]); 
    assign layer_0[8912] = in[19] ^ in[970]; 
    assign layer_0[8913] = in[465] | in[911]; 
    assign layer_0[8914] = ~in[257]; 
    assign layer_0[8915] = in[360] & ~in[618]; 
    assign layer_0[8916] = in[937]; 
    assign layer_0[8917] = ~in[84]; 
    assign layer_0[8918] = in[112] ^ in[365]; 
    assign layer_0[8919] = ~(in[503] | in[283]); 
    assign layer_0[8920] = in[906]; 
    assign layer_0[8921] = in[921]; 
    assign layer_0[8922] = in[299] & ~in[364]; 
    assign layer_0[8923] = in[715] & in[150]; 
    assign layer_0[8924] = ~(in[971] | in[63]); 
    assign layer_0[8925] = in[734] & ~in[177]; 
    assign layer_0[8926] = ~in[805] | (in[805] & in[286]); 
    assign layer_0[8927] = in[334] ^ in[844]; 
    assign layer_0[8928] = ~(in[50] | in[493]); 
    assign layer_0[8929] = ~(in[565] ^ in[843]); 
    assign layer_0[8930] = in[63]; 
    assign layer_0[8931] = in[663]; 
    assign layer_0[8932] = ~(in[463] ^ in[19]); 
    assign layer_0[8933] = in[809] ^ in[581]; 
    assign layer_0[8934] = in[589] ^ in[135]; 
    assign layer_0[8935] = ~in[1014]; 
    assign layer_0[8936] = ~(in[520] ^ in[804]); 
    assign layer_0[8937] = ~in[707]; 
    assign layer_0[8938] = in[711] ^ in[60]; 
    assign layer_0[8939] = ~in[396] | (in[656] & in[396]); 
    assign layer_0[8940] = ~(in[820] ^ in[933]); 
    assign layer_0[8941] = ~(in[350] ^ in[140]); 
    assign layer_0[8942] = ~in[492] | (in[281] & in[492]); 
    assign layer_0[8943] = ~(in[366] & in[616]); 
    assign layer_0[8944] = in[837]; 
    assign layer_0[8945] = in[750]; 
    assign layer_0[8946] = in[5] ^ in[250]; 
    assign layer_0[8947] = ~(in[570] ^ in[605]); 
    assign layer_0[8948] = in[805] & in[248]; 
    assign layer_0[8949] = in[441] ^ in[889]; 
    assign layer_0[8950] = ~in[166] | (in[166] & in[424]); 
    assign layer_0[8951] = ~(in[91] | in[315]); 
    assign layer_0[8952] = ~in[586]; 
    assign layer_0[8953] = ~(in[559] ^ in[705]); 
    assign layer_0[8954] = in[905] ^ in[899]; 
    assign layer_0[8955] = in[187] ^ in[1018]; 
    assign layer_0[8956] = in[540] & ~in[235]; 
    assign layer_0[8957] = in[789] | in[820]; 
    assign layer_0[8958] = in[357] | in[917]; 
    assign layer_0[8959] = ~in[266] | (in[266] & in[237]); 
    assign layer_0[8960] = in[759] & ~in[507]; 
    assign layer_0[8961] = ~in[1012] | (in[564] & in[1012]); 
    assign layer_0[8962] = ~in[727] | (in[727] & in[778]); 
    assign layer_0[8963] = ~(in[158] ^ in[13]); 
    assign layer_0[8964] = in[624] & in[138]; 
    assign layer_0[8965] = ~(in[602] ^ in[873]); 
    assign layer_0[8966] = ~(in[889] ^ in[858]); 
    assign layer_0[8967] = in[840] & ~in[834]; 
    assign layer_0[8968] = ~(in[724] ^ in[59]); 
    assign layer_0[8969] = ~(in[24] ^ in[576]); 
    assign layer_0[8970] = ~(in[348] ^ in[904]); 
    assign layer_0[8971] = ~(in[1015] ^ in[331]); 
    assign layer_0[8972] = in[747] ^ in[65]; 
    assign layer_0[8973] = in[456] ^ in[798]; 
    assign layer_0[8974] = in[522]; 
    assign layer_0[8975] = in[342] ^ in[829]; 
    assign layer_0[8976] = ~(in[948] ^ in[221]); 
    assign layer_0[8977] = ~(in[377] & in[309]); 
    assign layer_0[8978] = ~(in[563] ^ in[296]); 
    assign layer_0[8979] = in[51] & in[279]; 
    assign layer_0[8980] = ~(in[363] ^ in[566]); 
    assign layer_0[8981] = ~in[857] | (in[857] & in[144]); 
    assign layer_0[8982] = ~(in[243] ^ in[231]); 
    assign layer_0[8983] = in[488] ^ in[702]; 
    assign layer_0[8984] = in[264] ^ in[222]; 
    assign layer_0[8985] = ~(in[317] | in[823]); 
    assign layer_0[8986] = ~in[982] | (in[982] & in[1012]); 
    assign layer_0[8987] = ~in[163] | (in[576] & in[163]); 
    assign layer_0[8988] = in[323] ^ in[873]; 
    assign layer_0[8989] = ~in[599] | (in[599] & in[313]); 
    assign layer_0[8990] = 1'b1; 
    assign layer_0[8991] = in[598] ^ in[522]; 
    assign layer_0[8992] = in[548] & in[482]; 
    assign layer_0[8993] = in[966] | in[342]; 
    assign layer_0[8994] = in[654]; 
    assign layer_0[8995] = in[904]; 
    assign layer_0[8996] = ~(in[541] & in[748]); 
    assign layer_0[8997] = ~(in[448] | in[910]); 
    assign layer_0[8998] = in[703] ^ in[34]; 
    assign layer_0[8999] = in[379] | in[271]; 
    assign layer_0[9000] = ~(in[206] ^ in[623]); 
    assign layer_0[9001] = ~(in[524] ^ in[911]); 
    assign layer_0[9002] = in[422]; 
    assign layer_0[9003] = in[934] ^ in[857]; 
    assign layer_0[9004] = ~in[798] | (in[448] & in[798]); 
    assign layer_0[9005] = in[120]; 
    assign layer_0[9006] = in[1002]; 
    assign layer_0[9007] = ~in[922] | (in[922] & in[762]); 
    assign layer_0[9008] = ~in[240] | (in[240] & in[227]); 
    assign layer_0[9009] = ~(in[266] ^ in[29]); 
    assign layer_0[9010] = ~in[488] | (in[488] & in[243]); 
    assign layer_0[9011] = ~in[892]; 
    assign layer_0[9012] = ~in[195]; 
    assign layer_0[9013] = ~(in[612] | in[730]); 
    assign layer_0[9014] = ~(in[580] ^ in[34]); 
    assign layer_0[9015] = ~(in[811] | in[886]); 
    assign layer_0[9016] = ~in[730]; 
    assign layer_0[9017] = ~(in[280] ^ in[963]); 
    assign layer_0[9018] = in[284]; 
    assign layer_0[9019] = in[931]; 
    assign layer_0[9020] = in[81]; 
    assign layer_0[9021] = ~in[162] | (in[162] & in[948]); 
    assign layer_0[9022] = in[251] & in[482]; 
    assign layer_0[9023] = ~(in[775] ^ in[774]); 
    assign layer_0[9024] = ~in[691]; 
    assign layer_0[9025] = in[398] & ~in[247]; 
    assign layer_0[9026] = 1'b1; 
    assign layer_0[9027] = ~(in[823] ^ in[667]); 
    assign layer_0[9028] = ~(in[626] | in[987]); 
    assign layer_0[9029] = ~in[251] | (in[251] & in[485]); 
    assign layer_0[9030] = in[633]; 
    assign layer_0[9031] = ~(in[290] ^ in[144]); 
    assign layer_0[9032] = in[555] ^ in[936]; 
    assign layer_0[9033] = in[675]; 
    assign layer_0[9034] = in[583] ^ in[511]; 
    assign layer_0[9035] = ~(in[636] ^ in[221]); 
    assign layer_0[9036] = in[501] | in[267]; 
    assign layer_0[9037] = in[534] & ~in[524]; 
    assign layer_0[9038] = ~in[280] | (in[280] & in[937]); 
    assign layer_0[9039] = in[370] | in[599]; 
    assign layer_0[9040] = ~(in[951] ^ in[688]); 
    assign layer_0[9041] = in[319] | in[915]; 
    assign layer_0[9042] = in[6]; 
    assign layer_0[9043] = 1'b1; 
    assign layer_0[9044] = ~(in[91] | in[222]); 
    assign layer_0[9045] = in[157] & ~in[461]; 
    assign layer_0[9046] = ~(in[539] ^ in[354]); 
    assign layer_0[9047] = ~in[332] | (in[332] & in[13]); 
    assign layer_0[9048] = ~in[302] | (in[51] & in[302]); 
    assign layer_0[9049] = in[813] | in[477]; 
    assign layer_0[9050] = ~(in[949] ^ in[915]); 
    assign layer_0[9051] = in[723] | in[654]; 
    assign layer_0[9052] = in[101] & ~in[398]; 
    assign layer_0[9053] = ~(in[507] ^ in[142]); 
    assign layer_0[9054] = in[446]; 
    assign layer_0[9055] = in[76] & ~in[523]; 
    assign layer_0[9056] = ~(in[275] ^ in[261]); 
    assign layer_0[9057] = ~(in[807] ^ in[356]); 
    assign layer_0[9058] = in[706] ^ in[478]; 
    assign layer_0[9059] = ~in[842]; 
    assign layer_0[9060] = in[9] ^ in[1003]; 
    assign layer_0[9061] = in[476] ^ in[396]; 
    assign layer_0[9062] = in[856] ^ in[1001]; 
    assign layer_0[9063] = in[292] ^ in[877]; 
    assign layer_0[9064] = in[163] & ~in[302]; 
    assign layer_0[9065] = ~(in[99] ^ in[29]); 
    assign layer_0[9066] = ~(in[66] | in[961]); 
    assign layer_0[9067] = ~in[422] | (in[966] & in[422]); 
    assign layer_0[9068] = in[147] ^ in[216]; 
    assign layer_0[9069] = ~(in[919] ^ in[886]); 
    assign layer_0[9070] = in[254] ^ in[74]; 
    assign layer_0[9071] = in[827] ^ in[923]; 
    assign layer_0[9072] = ~in[539]; 
    assign layer_0[9073] = ~(in[386] ^ in[902]); 
    assign layer_0[9074] = ~in[899]; 
    assign layer_0[9075] = in[761] ^ in[824]; 
    assign layer_0[9076] = in[669] & ~in[233]; 
    assign layer_0[9077] = in[951] & in[410]; 
    assign layer_0[9078] = in[98] | in[35]; 
    assign layer_0[9079] = ~in[397] | (in[262] & in[397]); 
    assign layer_0[9080] = in[838] | in[162]; 
    assign layer_0[9081] = in[129] ^ in[935]; 
    assign layer_0[9082] = in[44] | in[985]; 
    assign layer_0[9083] = ~in[488] | (in[488] & in[606]); 
    assign layer_0[9084] = ~(in[677] ^ in[311]); 
    assign layer_0[9085] = in[598] | in[3]; 
    assign layer_0[9086] = ~in[724]; 
    assign layer_0[9087] = ~in[1000] | (in[530] & in[1000]); 
    assign layer_0[9088] = in[882] | in[929]; 
    assign layer_0[9089] = in[275] ^ in[1015]; 
    assign layer_0[9090] = in[925] ^ in[795]; 
    assign layer_0[9091] = ~(in[317] ^ in[509]); 
    assign layer_0[9092] = in[679] & in[645]; 
    assign layer_0[9093] = ~(in[625] ^ in[541]); 
    assign layer_0[9094] = in[365] | in[154]; 
    assign layer_0[9095] = ~(in[811] ^ in[734]); 
    assign layer_0[9096] = ~in[159] | (in[159] & in[239]); 
    assign layer_0[9097] = ~(in[82] ^ in[762]); 
    assign layer_0[9098] = ~(in[822] & in[932]); 
    assign layer_0[9099] = in[476] & ~in[931]; 
    assign layer_0[9100] = in[415] & ~in[985]; 
    assign layer_0[9101] = in[251] & in[228]; 
    assign layer_0[9102] = in[319] ^ in[342]; 
    assign layer_0[9103] = in[758] & ~in[436]; 
    assign layer_0[9104] = in[779] | in[311]; 
    assign layer_0[9105] = in[359] ^ in[8]; 
    assign layer_0[9106] = ~in[24] | (in[24] & in[522]); 
    assign layer_0[9107] = in[156] & ~in[141]; 
    assign layer_0[9108] = ~(in[513] ^ in[952]); 
    assign layer_0[9109] = 1'b1; 
    assign layer_0[9110] = ~in[326]; 
    assign layer_0[9111] = in[921] ^ in[962]; 
    assign layer_0[9112] = ~(in[215] & in[396]); 
    assign layer_0[9113] = ~in[745] | (in[745] & in[12]); 
    assign layer_0[9114] = in[249] & ~in[935]; 
    assign layer_0[9115] = ~(in[1013] ^ in[756]); 
    assign layer_0[9116] = ~(in[694] ^ in[493]); 
    assign layer_0[9117] = in[874] & in[795]; 
    assign layer_0[9118] = in[431] & in[407]; 
    assign layer_0[9119] = ~(in[711] & in[613]); 
    assign layer_0[9120] = ~(in[729] ^ in[732]); 
    assign layer_0[9121] = ~(in[859] ^ in[498]); 
    assign layer_0[9122] = ~in[600]; 
    assign layer_0[9123] = 1'b0; 
    assign layer_0[9124] = in[789] & in[121]; 
    assign layer_0[9125] = in[123] ^ in[934]; 
    assign layer_0[9126] = in[566] ^ in[381]; 
    assign layer_0[9127] = 1'b1; 
    assign layer_0[9128] = in[963] | in[574]; 
    assign layer_0[9129] = ~in[119] | (in[119] & in[218]); 
    assign layer_0[9130] = ~in[801]; 
    assign layer_0[9131] = ~in[893] | (in[30] & in[893]); 
    assign layer_0[9132] = ~in[967] | (in[790] & in[967]); 
    assign layer_0[9133] = in[655] ^ in[631]; 
    assign layer_0[9134] = ~in[138]; 
    assign layer_0[9135] = in[409] & ~in[627]; 
    assign layer_0[9136] = in[1017] ^ in[730]; 
    assign layer_0[9137] = ~(in[757] ^ in[378]); 
    assign layer_0[9138] = ~(in[937] ^ in[965]); 
    assign layer_0[9139] = in[1017] ^ in[793]; 
    assign layer_0[9140] = ~in[837]; 
    assign layer_0[9141] = in[891]; 
    assign layer_0[9142] = ~in[222]; 
    assign layer_0[9143] = ~(in[925] & in[667]); 
    assign layer_0[9144] = in[423] & ~in[911]; 
    assign layer_0[9145] = ~in[894]; 
    assign layer_0[9146] = ~(in[886] ^ in[888]); 
    assign layer_0[9147] = in[986]; 
    assign layer_0[9148] = in[295]; 
    assign layer_0[9149] = ~in[243]; 
    assign layer_0[9150] = in[884] ^ in[587]; 
    assign layer_0[9151] = ~in[223]; 
    assign layer_0[9152] = 1'b1; 
    assign layer_0[9153] = in[595] & ~in[672]; 
    assign layer_0[9154] = ~(in[882] ^ in[1002]); 
    assign layer_0[9155] = ~(in[616] & in[348]); 
    assign layer_0[9156] = ~(in[892] | in[995]); 
    assign layer_0[9157] = in[521] ^ in[807]; 
    assign layer_0[9158] = ~(in[904] | in[266]); 
    assign layer_0[9159] = ~(in[650] | in[819]); 
    assign layer_0[9160] = in[678] & ~in[429]; 
    assign layer_0[9161] = in[629] ^ in[597]; 
    assign layer_0[9162] = in[549] & in[275]; 
    assign layer_0[9163] = in[838] ^ in[855]; 
    assign layer_0[9164] = ~(in[758] ^ in[460]); 
    assign layer_0[9165] = ~(in[633] & in[586]); 
    assign layer_0[9166] = ~(in[905] | in[547]); 
    assign layer_0[9167] = in[418] ^ in[49]; 
    assign layer_0[9168] = ~(in[387] | in[416]); 
    assign layer_0[9169] = ~in[77] | (in[879] & in[77]); 
    assign layer_0[9170] = in[38]; 
    assign layer_0[9171] = ~(in[17] | in[353]); 
    assign layer_0[9172] = in[714] & in[523]; 
    assign layer_0[9173] = in[958] ^ in[910]; 
    assign layer_0[9174] = ~in[623]; 
    assign layer_0[9175] = ~(in[723] ^ in[808]); 
    assign layer_0[9176] = in[875]; 
    assign layer_0[9177] = in[823] & ~in[837]; 
    assign layer_0[9178] = in[109] ^ in[591]; 
    assign layer_0[9179] = ~in[285]; 
    assign layer_0[9180] = ~in[969]; 
    assign layer_0[9181] = in[596]; 
    assign layer_0[9182] = in[1018]; 
    assign layer_0[9183] = ~(in[808] ^ in[825]); 
    assign layer_0[9184] = ~(in[631] ^ in[899]); 
    assign layer_0[9185] = ~(in[263] ^ in[645]); 
    assign layer_0[9186] = ~in[444]; 
    assign layer_0[9187] = ~in[477]; 
    assign layer_0[9188] = ~(in[657] ^ in[601]); 
    assign layer_0[9189] = ~(in[889] | in[522]); 
    assign layer_0[9190] = in[602] | in[555]; 
    assign layer_0[9191] = in[837] ^ in[257]; 
    assign layer_0[9192] = in[891] & ~in[873]; 
    assign layer_0[9193] = 1'b1; 
    assign layer_0[9194] = in[264] & in[973]; 
    assign layer_0[9195] = in[966]; 
    assign layer_0[9196] = ~in[404]; 
    assign layer_0[9197] = in[800] | in[888]; 
    assign layer_0[9198] = in[803] | in[952]; 
    assign layer_0[9199] = in[340] ^ in[420]; 
    assign layer_0[9200] = in[242] | in[329]; 
    assign layer_0[9201] = ~(in[429] | in[901]); 
    assign layer_0[9202] = in[534]; 
    assign layer_0[9203] = in[694] & ~in[521]; 
    assign layer_0[9204] = in[857] & ~in[559]; 
    assign layer_0[9205] = in[369] | in[312]; 
    assign layer_0[9206] = in[264]; 
    assign layer_0[9207] = in[734] & ~in[959]; 
    assign layer_0[9208] = ~in[723] | (in[723] & in[487]); 
    assign layer_0[9209] = in[603] | in[708]; 
    assign layer_0[9210] = ~in[352] | (in[675] & in[352]); 
    assign layer_0[9211] = ~(in[470] | in[840]); 
    assign layer_0[9212] = in[296] & ~in[208]; 
    assign layer_0[9213] = in[570] & ~in[640]; 
    assign layer_0[9214] = in[646] & ~in[331]; 
    assign layer_0[9215] = ~in[722] | (in[722] & in[21]); 
    assign layer_0[9216] = ~(in[406] ^ in[844]); 
    assign layer_0[9217] = in[996] | in[757]; 
    assign layer_0[9218] = ~in[948]; 
    assign layer_0[9219] = ~(in[129] ^ in[970]); 
    assign layer_0[9220] = in[724] | in[967]; 
    assign layer_0[9221] = ~(in[475] & in[383]); 
    assign layer_0[9222] = in[324] | in[877]; 
    assign layer_0[9223] = in[685] | in[594]; 
    assign layer_0[9224] = ~in[146]; 
    assign layer_0[9225] = ~in[155]; 
    assign layer_0[9226] = ~in[642]; 
    assign layer_0[9227] = in[690] ^ in[868]; 
    assign layer_0[9228] = ~in[594]; 
    assign layer_0[9229] = in[572] & ~in[762]; 
    assign layer_0[9230] = ~(in[622] & in[131]); 
    assign layer_0[9231] = in[583] | in[491]; 
    assign layer_0[9232] = ~(in[877] | in[553]); 
    assign layer_0[9233] = ~in[807]; 
    assign layer_0[9234] = ~(in[266] ^ in[825]); 
    assign layer_0[9235] = ~(in[1019] | in[613]); 
    assign layer_0[9236] = ~in[466] | (in[1004] & in[466]); 
    assign layer_0[9237] = ~in[885]; 
    assign layer_0[9238] = in[539] ^ in[700]; 
    assign layer_0[9239] = in[788] & in[437]; 
    assign layer_0[9240] = in[810] | in[733]; 
    assign layer_0[9241] = in[421] & in[554]; 
    assign layer_0[9242] = in[884] ^ in[939]; 
    assign layer_0[9243] = ~in[976] | (in[976] & in[765]); 
    assign layer_0[9244] = in[175] & in[240]; 
    assign layer_0[9245] = ~(in[939] ^ in[63]); 
    assign layer_0[9246] = in[552] & ~in[430]; 
    assign layer_0[9247] = in[502] & in[50]; 
    assign layer_0[9248] = in[18] | in[382]; 
    assign layer_0[9249] = in[759] ^ in[509]; 
    assign layer_0[9250] = in[56] ^ in[30]; 
    assign layer_0[9251] = ~(in[662] ^ in[382]); 
    assign layer_0[9252] = ~in[886] | (in[160] & in[886]); 
    assign layer_0[9253] = ~in[667] | (in[520] & in[667]); 
    assign layer_0[9254] = ~(in[85] ^ in[941]); 
    assign layer_0[9255] = ~(in[852] | in[62]); 
    assign layer_0[9256] = in[230] & ~in[252]; 
    assign layer_0[9257] = ~(in[450] & in[202]); 
    assign layer_0[9258] = in[61] ^ in[759]; 
    assign layer_0[9259] = ~(in[665] ^ in[261]); 
    assign layer_0[9260] = ~(in[983] | in[805]); 
    assign layer_0[9261] = ~(in[939] ^ in[890]); 
    assign layer_0[9262] = in[952] ^ in[920]; 
    assign layer_0[9263] = in[739] | in[509]; 
    assign layer_0[9264] = in[287]; 
    assign layer_0[9265] = ~in[887] | (in[887] & in[493]); 
    assign layer_0[9266] = in[707] | in[448]; 
    assign layer_0[9267] = in[619] & ~in[331]; 
    assign layer_0[9268] = in[28] & in[310]; 
    assign layer_0[9269] = in[517] ^ in[296]; 
    assign layer_0[9270] = in[985] & in[454]; 
    assign layer_0[9271] = ~in[777] | (in[922] & in[777]); 
    assign layer_0[9272] = ~(in[620] ^ in[1004]); 
    assign layer_0[9273] = in[668]; 
    assign layer_0[9274] = in[924] & ~in[959]; 
    assign layer_0[9275] = in[109] ^ in[493]; 
    assign layer_0[9276] = ~in[853] | (in[234] & in[853]); 
    assign layer_0[9277] = ~(in[1022] | in[207]); 
    assign layer_0[9278] = ~(in[699] & in[245]); 
    assign layer_0[9279] = in[229] ^ in[262]; 
    assign layer_0[9280] = ~in[4] | (in[4] & in[667]); 
    assign layer_0[9281] = ~(in[724] ^ in[147]); 
    assign layer_0[9282] = in[603] | in[722]; 
    assign layer_0[9283] = in[982] & in[824]; 
    assign layer_0[9284] = in[493] & in[482]; 
    assign layer_0[9285] = ~(in[757] | in[772]); 
    assign layer_0[9286] = in[889] | in[580]; 
    assign layer_0[9287] = ~(in[198] | in[989]); 
    assign layer_0[9288] = in[829] | in[659]; 
    assign layer_0[9289] = in[518] ^ in[413]; 
    assign layer_0[9290] = in[948] ^ in[935]; 
    assign layer_0[9291] = ~(in[239] | in[1018]); 
    assign layer_0[9292] = ~(in[251] ^ in[148]); 
    assign layer_0[9293] = in[839]; 
    assign layer_0[9294] = ~in[201] | (in[201] & in[14]); 
    assign layer_0[9295] = ~(in[667] | in[902]); 
    assign layer_0[9296] = ~(in[937] ^ in[648]); 
    assign layer_0[9297] = ~in[62] | (in[62] & in[322]); 
    assign layer_0[9298] = ~(in[296] ^ in[262]); 
    assign layer_0[9299] = ~in[935]; 
    assign layer_0[9300] = ~(in[573] | in[575]); 
    assign layer_0[9301] = in[728]; 
    assign layer_0[9302] = ~in[219] | (in[522] & in[219]); 
    assign layer_0[9303] = in[159] & ~in[872]; 
    assign layer_0[9304] = ~in[78]; 
    assign layer_0[9305] = in[225] ^ in[355]; 
    assign layer_0[9306] = 1'b0; 
    assign layer_0[9307] = ~(in[628] ^ in[689]); 
    assign layer_0[9308] = ~(in[491] | in[1003]); 
    assign layer_0[9309] = ~in[632] | (in[819] & in[632]); 
    assign layer_0[9310] = ~(in[45] ^ in[375]); 
    assign layer_0[9311] = in[761] ^ in[999]; 
    assign layer_0[9312] = in[390] & ~in[977]; 
    assign layer_0[9313] = ~(in[732] ^ in[602]); 
    assign layer_0[9314] = ~(in[597] ^ in[907]); 
    assign layer_0[9315] = ~(in[859] | in[463]); 
    assign layer_0[9316] = in[299]; 
    assign layer_0[9317] = ~in[505] | (in[495] & in[505]); 
    assign layer_0[9318] = ~in[691] | (in[691] & in[323]); 
    assign layer_0[9319] = in[915] ^ in[953]; 
    assign layer_0[9320] = in[524] ^ in[507]; 
    assign layer_0[9321] = in[908] & ~in[743]; 
    assign layer_0[9322] = in[501] & ~in[110]; 
    assign layer_0[9323] = in[45] | in[141]; 
    assign layer_0[9324] = in[858] & in[857]; 
    assign layer_0[9325] = ~(in[324] ^ in[1016]); 
    assign layer_0[9326] = in[611] ^ in[869]; 
    assign layer_0[9327] = in[318] ^ in[952]; 
    assign layer_0[9328] = in[727] & ~in[822]; 
    assign layer_0[9329] = 1'b0; 
    assign layer_0[9330] = ~(in[11] ^ in[693]); 
    assign layer_0[9331] = ~(in[597] ^ in[963]); 
    assign layer_0[9332] = ~in[689] | (in[900] & in[689]); 
    assign layer_0[9333] = ~(in[85] ^ in[73]); 
    assign layer_0[9334] = in[743] ^ in[887]; 
    assign layer_0[9335] = ~in[638] | (in[638] & in[611]); 
    assign layer_0[9336] = ~(in[862] | in[943]); 
    assign layer_0[9337] = ~(in[615] ^ in[616]); 
    assign layer_0[9338] = in[252] ^ in[662]; 
    assign layer_0[9339] = in[760] & ~in[985]; 
    assign layer_0[9340] = ~(in[980] | in[473]); 
    assign layer_0[9341] = in[18] ^ in[445]; 
    assign layer_0[9342] = ~in[854]; 
    assign layer_0[9343] = ~(in[508] ^ in[254]); 
    assign layer_0[9344] = ~in[819]; 
    assign layer_0[9345] = in[436]; 
    assign layer_0[9346] = ~in[338]; 
    assign layer_0[9347] = in[649] ^ in[743]; 
    assign layer_0[9348] = ~(in[740] & in[451]); 
    assign layer_0[9349] = in[36] & in[517]; 
    assign layer_0[9350] = in[998] & in[969]; 
    assign layer_0[9351] = ~(in[869] ^ in[519]); 
    assign layer_0[9352] = ~in[188]; 
    assign layer_0[9353] = ~(in[721] ^ in[611]); 
    assign layer_0[9354] = in[218] ^ in[613]; 
    assign layer_0[9355] = in[332] & ~in[780]; 
    assign layer_0[9356] = in[95] & ~in[84]; 
    assign layer_0[9357] = in[1001] & ~in[303]; 
    assign layer_0[9358] = ~(in[917] ^ in[903]); 
    assign layer_0[9359] = ~(in[952] ^ in[955]); 
    assign layer_0[9360] = ~(in[78] ^ in[126]); 
    assign layer_0[9361] = ~(in[548] ^ in[867]); 
    assign layer_0[9362] = ~(in[599] ^ in[319]); 
    assign layer_0[9363] = in[683] & in[657]; 
    assign layer_0[9364] = 1'b0; 
    assign layer_0[9365] = in[842] ^ in[699]; 
    assign layer_0[9366] = in[859] ^ in[158]; 
    assign layer_0[9367] = in[854] ^ in[676]; 
    assign layer_0[9368] = ~(in[165] ^ in[894]); 
    assign layer_0[9369] = ~(in[921] ^ in[715]); 
    assign layer_0[9370] = in[823] | in[667]; 
    assign layer_0[9371] = in[835]; 
    assign layer_0[9372] = in[366]; 
    assign layer_0[9373] = in[557] ^ in[147]; 
    assign layer_0[9374] = ~(in[665] ^ in[396]); 
    assign layer_0[9375] = in[728] & ~in[514]; 
    assign layer_0[9376] = in[602] ^ in[579]; 
    assign layer_0[9377] = in[64] ^ in[744]; 
    assign layer_0[9378] = in[961] ^ in[312]; 
    assign layer_0[9379] = in[28] & ~in[854]; 
    assign layer_0[9380] = ~in[729] | (in[339] & in[729]); 
    assign layer_0[9381] = ~in[209]; 
    assign layer_0[9382] = in[173] & in[569]; 
    assign layer_0[9383] = in[592] & in[55]; 
    assign layer_0[9384] = in[438]; 
    assign layer_0[9385] = in[639]; 
    assign layer_0[9386] = ~in[906] | (in[906] & in[898]); 
    assign layer_0[9387] = in[717]; 
    assign layer_0[9388] = ~(in[413] ^ in[406]); 
    assign layer_0[9389] = ~in[952] | (in[952] & in[547]); 
    assign layer_0[9390] = ~(in[413] | in[1017]); 
    assign layer_0[9391] = in[12] ^ in[248]; 
    assign layer_0[9392] = in[674] ^ in[708]; 
    assign layer_0[9393] = in[223] & ~in[846]; 
    assign layer_0[9394] = ~(in[919] & in[711]); 
    assign layer_0[9395] = ~(in[555] ^ in[652]); 
    assign layer_0[9396] = in[604] & ~in[260]; 
    assign layer_0[9397] = in[572] ^ in[620]; 
    assign layer_0[9398] = in[633] & ~in[713]; 
    assign layer_0[9399] = ~in[993] | (in[666] & in[993]); 
    assign layer_0[9400] = in[94] ^ in[931]; 
    assign layer_0[9401] = ~in[371] | (in[371] & in[174]); 
    assign layer_0[9402] = in[870] ^ in[951]; 
    assign layer_0[9403] = in[224]; 
    assign layer_0[9404] = in[79] ^ in[529]; 
    assign layer_0[9405] = ~in[598] | (in[915] & in[598]); 
    assign layer_0[9406] = ~(in[16] | in[215]); 
    assign layer_0[9407] = in[125] & ~in[809]; 
    assign layer_0[9408] = ~(in[874] ^ in[603]); 
    assign layer_0[9409] = in[84] & ~in[461]; 
    assign layer_0[9410] = ~(in[610] & in[237]); 
    assign layer_0[9411] = in[872] ^ in[502]; 
    assign layer_0[9412] = ~in[29] | (in[883] & in[29]); 
    assign layer_0[9413] = ~in[690] | (in[690] & in[554]); 
    assign layer_0[9414] = ~(in[615] ^ in[749]); 
    assign layer_0[9415] = in[899] ^ in[518]; 
    assign layer_0[9416] = in[142] ^ in[283]; 
    assign layer_0[9417] = ~in[607] | (in[885] & in[607]); 
    assign layer_0[9418] = ~(in[259] ^ in[253]); 
    assign layer_0[9419] = ~(in[341] ^ in[734]); 
    assign layer_0[9420] = in[317] ^ in[51]; 
    assign layer_0[9421] = in[483] & ~in[303]; 
    assign layer_0[9422] = ~in[264] | (in[30] & in[264]); 
    assign layer_0[9423] = ~(in[344] ^ in[949]); 
    assign layer_0[9424] = ~(in[357] ^ in[216]); 
    assign layer_0[9425] = in[926]; 
    assign layer_0[9426] = ~(in[876] & in[576]); 
    assign layer_0[9427] = ~(in[573] ^ in[840]); 
    assign layer_0[9428] = in[761] & in[761]; 
    assign layer_0[9429] = ~in[977] | (in[977] & in[546]); 
    assign layer_0[9430] = ~(in[731] & in[775]); 
    assign layer_0[9431] = in[597] ^ in[485]; 
    assign layer_0[9432] = in[341] | in[882]; 
    assign layer_0[9433] = ~(in[792] | in[831]); 
    assign layer_0[9434] = ~(in[836] ^ in[842]); 
    assign layer_0[9435] = in[708]; 
    assign layer_0[9436] = ~in[537] | (in[537] & in[354]); 
    assign layer_0[9437] = ~in[614]; 
    assign layer_0[9438] = ~in[874] | (in[874] & in[347]); 
    assign layer_0[9439] = in[1004] | in[622]; 
    assign layer_0[9440] = in[165] & ~in[74]; 
    assign layer_0[9441] = in[721] ^ in[562]; 
    assign layer_0[9442] = in[245] & ~in[627]; 
    assign layer_0[9443] = ~(in[659] ^ in[436]); 
    assign layer_0[9444] = in[353] & in[112]; 
    assign layer_0[9445] = in[254]; 
    assign layer_0[9446] = in[444] ^ in[4]; 
    assign layer_0[9447] = in[947]; 
    assign layer_0[9448] = ~(in[749] ^ in[322]); 
    assign layer_0[9449] = in[782] & ~in[816]; 
    assign layer_0[9450] = 1'b0; 
    assign layer_0[9451] = ~(in[708] ^ in[237]); 
    assign layer_0[9452] = in[503] ^ in[499]; 
    assign layer_0[9453] = 1'b0; 
    assign layer_0[9454] = ~(in[60] & in[114]); 
    assign layer_0[9455] = ~(in[322] ^ in[646]); 
    assign layer_0[9456] = ~in[468]; 
    assign layer_0[9457] = in[355] ^ in[583]; 
    assign layer_0[9458] = ~(in[954] ^ in[904]); 
    assign layer_0[9459] = in[192] & in[310]; 
    assign layer_0[9460] = ~(in[997] | in[980]); 
    assign layer_0[9461] = ~(in[764] ^ in[713]); 
    assign layer_0[9462] = ~(in[418] ^ in[955]); 
    assign layer_0[9463] = in[335] ^ in[730]; 
    assign layer_0[9464] = in[669] | in[210]; 
    assign layer_0[9465] = ~in[501] | (in[62] & in[501]); 
    assign layer_0[9466] = ~(in[997] ^ in[290]); 
    assign layer_0[9467] = ~(in[564] ^ in[838]); 
    assign layer_0[9468] = in[172] ^ in[354]; 
    assign layer_0[9469] = ~(in[232] & in[332]); 
    assign layer_0[9470] = ~(in[739] | in[612]); 
    assign layer_0[9471] = ~(in[715] ^ in[775]); 
    assign layer_0[9472] = in[504] & in[379]; 
    assign layer_0[9473] = in[520] ^ in[835]; 
    assign layer_0[9474] = ~(in[692] | in[643]); 
    assign layer_0[9475] = ~(in[964] ^ in[602]); 
    assign layer_0[9476] = ~(in[776] ^ in[75]); 
    assign layer_0[9477] = in[582] & ~in[1010]; 
    assign layer_0[9478] = in[708] ^ in[715]; 
    assign layer_0[9479] = ~(in[306] ^ in[327]); 
    assign layer_0[9480] = ~in[613]; 
    assign layer_0[9481] = ~in[248]; 
    assign layer_0[9482] = ~in[260] | (in[873] & in[260]); 
    assign layer_0[9483] = in[1007] ^ in[510]; 
    assign layer_0[9484] = ~(in[838] | in[867]); 
    assign layer_0[9485] = in[504] & ~in[691]; 
    assign layer_0[9486] = in[132]; 
    assign layer_0[9487] = in[934] ^ in[547]; 
    assign layer_0[9488] = ~(in[266] ^ in[729]); 
    assign layer_0[9489] = in[381] ^ in[63]; 
    assign layer_0[9490] = in[231] | in[330]; 
    assign layer_0[9491] = in[859] ^ in[886]; 
    assign layer_0[9492] = ~in[320]; 
    assign layer_0[9493] = ~(in[233] ^ in[820]); 
    assign layer_0[9494] = in[773] ^ in[742]; 
    assign layer_0[9495] = ~(in[691] ^ in[679]); 
    assign layer_0[9496] = ~(in[704] & in[495]); 
    assign layer_0[9497] = in[872] | in[867]; 
    assign layer_0[9498] = in[584] | in[284]; 
    assign layer_0[9499] = in[411] ^ in[207]; 
    assign layer_0[9500] = ~(in[776] | in[656]); 
    assign layer_0[9501] = in[656] ^ in[310]; 
    assign layer_0[9502] = in[110]; 
    assign layer_0[9503] = ~in[696] | (in[696] & in[34]); 
    assign layer_0[9504] = in[517]; 
    assign layer_0[9505] = ~in[190]; 
    assign layer_0[9506] = in[479] | in[652]; 
    assign layer_0[9507] = ~(in[584] ^ in[874]); 
    assign layer_0[9508] = ~(in[341] & in[663]); 
    assign layer_0[9509] = in[182] & ~in[1000]; 
    assign layer_0[9510] = in[270] ^ in[210]; 
    assign layer_0[9511] = in[655] ^ in[894]; 
    assign layer_0[9512] = in[880] | in[339]; 
    assign layer_0[9513] = in[603]; 
    assign layer_0[9514] = ~in[477] | (in[167] & in[477]); 
    assign layer_0[9515] = ~(in[839] ^ in[500]); 
    assign layer_0[9516] = ~in[368] | (in[491] & in[368]); 
    assign layer_0[9517] = ~in[676] | (in[334] & in[676]); 
    assign layer_0[9518] = ~(in[969] ^ in[262]); 
    assign layer_0[9519] = in[252] & in[338]; 
    assign layer_0[9520] = in[894] ^ in[910]; 
    assign layer_0[9521] = in[173] ^ in[163]; 
    assign layer_0[9522] = ~(in[820] ^ in[241]); 
    assign layer_0[9523] = ~(in[482] & in[407]); 
    assign layer_0[9524] = ~(in[613] ^ in[618]); 
    assign layer_0[9525] = in[641] & in[345]; 
    assign layer_0[9526] = ~in[24] | (in[24] & in[754]); 
    assign layer_0[9527] = in[119] & ~in[958]; 
    assign layer_0[9528] = ~in[156] | (in[156] & in[78]); 
    assign layer_0[9529] = in[540] | in[349]; 
    assign layer_0[9530] = 1'b1; 
    assign layer_0[9531] = ~in[653] | (in[653] & in[354]); 
    assign layer_0[9532] = in[538] ^ in[300]; 
    assign layer_0[9533] = ~(in[570] ^ in[714]); 
    assign layer_0[9534] = ~(in[921] ^ in[668]); 
    assign layer_0[9535] = in[724] ^ in[67]; 
    assign layer_0[9536] = ~(in[699] ^ in[941]); 
    assign layer_0[9537] = ~in[1017]; 
    assign layer_0[9538] = in[800] ^ in[745]; 
    assign layer_0[9539] = ~(in[247] & in[10]); 
    assign layer_0[9540] = ~in[1016] | (in[1016] & in[719]); 
    assign layer_0[9541] = ~in[519] | (in[922] & in[519]); 
    assign layer_0[9542] = 1'b1; 
    assign layer_0[9543] = in[808] ^ in[500]; 
    assign layer_0[9544] = ~(in[905] ^ in[903]); 
    assign layer_0[9545] = ~in[291]; 
    assign layer_0[9546] = in[114]; 
    assign layer_0[9547] = in[534] ^ in[410]; 
    assign layer_0[9548] = ~in[581] | (in[581] & in[239]); 
    assign layer_0[9549] = in[948] ^ in[311]; 
    assign layer_0[9550] = in[187]; 
    assign layer_0[9551] = ~in[176]; 
    assign layer_0[9552] = ~(in[684] ^ in[317]); 
    assign layer_0[9553] = ~in[953] | (in[659] & in[953]); 
    assign layer_0[9554] = ~in[818] | (in[818] & in[425]); 
    assign layer_0[9555] = in[910] ^ in[897]; 
    assign layer_0[9556] = in[455] & in[638]; 
    assign layer_0[9557] = ~in[711] | (in[711] & in[333]); 
    assign layer_0[9558] = in[612]; 
    assign layer_0[9559] = ~(in[726] ^ in[869]); 
    assign layer_0[9560] = ~(in[644] & in[580]); 
    assign layer_0[9561] = in[476] & in[549]; 
    assign layer_0[9562] = ~(in[776] | in[793]); 
    assign layer_0[9563] = ~(in[937] ^ in[936]); 
    assign layer_0[9564] = in[491] & ~in[965]; 
    assign layer_0[9565] = ~(in[741] ^ in[78]); 
    assign layer_0[9566] = ~(in[810] ^ in[728]); 
    assign layer_0[9567] = ~(in[333] ^ in[934]); 
    assign layer_0[9568] = ~in[373]; 
    assign layer_0[9569] = ~in[917]; 
    assign layer_0[9570] = ~(in[886] ^ in[878]); 
    assign layer_0[9571] = in[98] & ~in[873]; 
    assign layer_0[9572] = ~in[876] | (in[502] & in[876]); 
    assign layer_0[9573] = ~(in[471] ^ in[722]); 
    assign layer_0[9574] = in[766] | in[484]; 
    assign layer_0[9575] = ~(in[982] ^ in[243]); 
    assign layer_0[9576] = ~in[503]; 
    assign layer_0[9577] = 1'b0; 
    assign layer_0[9578] = in[118] & in[978]; 
    assign layer_0[9579] = in[226] ^ in[130]; 
    assign layer_0[9580] = ~(in[698] | in[287]); 
    assign layer_0[9581] = in[930] ^ in[672]; 
    assign layer_0[9582] = in[738] & in[465]; 
    assign layer_0[9583] = in[827] ^ in[808]; 
    assign layer_0[9584] = ~(in[664] ^ in[492]); 
    assign layer_0[9585] = ~(in[704] ^ in[586]); 
    assign layer_0[9586] = in[714] ^ in[712]; 
    assign layer_0[9587] = ~(in[614] ^ in[236]); 
    assign layer_0[9588] = ~(in[205] ^ in[222]); 
    assign layer_0[9589] = in[675] & ~in[341]; 
    assign layer_0[9590] = in[910] & ~in[771]; 
    assign layer_0[9591] = ~(in[960] | in[352]); 
    assign layer_0[9592] = in[299] ^ in[705]; 
    assign layer_0[9593] = ~in[83]; 
    assign layer_0[9594] = ~in[108]; 
    assign layer_0[9595] = in[269] ^ in[181]; 
    assign layer_0[9596] = ~(in[710] ^ in[203]); 
    assign layer_0[9597] = ~(in[851] | in[985]); 
    assign layer_0[9598] = in[921] ^ in[903]; 
    assign layer_0[9599] = ~(in[873] | in[717]); 
    assign layer_0[9600] = in[361] & in[586]; 
    assign layer_0[9601] = ~in[951] | (in[951] & in[762]); 
    assign layer_0[9602] = ~in[436] | (in[843] & in[436]); 
    assign layer_0[9603] = ~(in[792] & in[806]); 
    assign layer_0[9604] = ~in[868] | (in[319] & in[868]); 
    assign layer_0[9605] = in[604] & in[312]; 
    assign layer_0[9606] = ~(in[755] | in[18]); 
    assign layer_0[9607] = in[175] ^ in[382]; 
    assign layer_0[9608] = in[889]; 
    assign layer_0[9609] = in[698]; 
    assign layer_0[9610] = ~in[968] | (in[968] & in[860]); 
    assign layer_0[9611] = in[253] ^ in[943]; 
    assign layer_0[9612] = ~(in[606] | in[77]); 
    assign layer_0[9613] = in[440] & ~in[192]; 
    assign layer_0[9614] = in[536] & in[853]; 
    assign layer_0[9615] = ~(in[138] | in[141]); 
    assign layer_0[9616] = ~(in[460] ^ in[616]); 
    assign layer_0[9617] = in[267] ^ in[82]; 
    assign layer_0[9618] = ~in[330] | (in[330] & in[375]); 
    assign layer_0[9619] = in[588] ^ in[710]; 
    assign layer_0[9620] = ~in[756] | (in[756] & in[159]); 
    assign layer_0[9621] = ~in[995]; 
    assign layer_0[9622] = ~in[313] | (in[550] & in[313]); 
    assign layer_0[9623] = ~in[29]; 
    assign layer_0[9624] = ~in[780]; 
    assign layer_0[9625] = in[708]; 
    assign layer_0[9626] = in[636] & in[446]; 
    assign layer_0[9627] = ~in[379]; 
    assign layer_0[9628] = ~in[317] | (in[317] & in[730]); 
    assign layer_0[9629] = ~in[836]; 
    assign layer_0[9630] = in[808] | in[809]; 
    assign layer_0[9631] = in[732]; 
    assign layer_0[9632] = ~(in[41] ^ in[607]); 
    assign layer_0[9633] = in[966] ^ in[807]; 
    assign layer_0[9634] = ~(in[628] ^ in[653]); 
    assign layer_0[9635] = in[708] & ~in[754]; 
    assign layer_0[9636] = ~(in[739] ^ in[4]); 
    assign layer_0[9637] = in[972] | in[943]; 
    assign layer_0[9638] = ~(in[253] ^ in[603]); 
    assign layer_0[9639] = in[455] & in[103]; 
    assign layer_0[9640] = in[633]; 
    assign layer_0[9641] = in[999] ^ in[983]; 
    assign layer_0[9642] = in[473]; 
    assign layer_0[9643] = ~in[900]; 
    assign layer_0[9644] = in[512] & ~in[157]; 
    assign layer_0[9645] = in[36]; 
    assign layer_0[9646] = ~(in[660] & in[503]); 
    assign layer_0[9647] = ~in[580]; 
    assign layer_0[9648] = ~(in[563] | in[625]); 
    assign layer_0[9649] = in[160] & ~in[595]; 
    assign layer_0[9650] = in[647] ^ in[145]; 
    assign layer_0[9651] = ~in[874]; 
    assign layer_0[9652] = ~in[504] | (in[504] & in[779]); 
    assign layer_0[9653] = ~in[176] | (in[643] & in[176]); 
    assign layer_0[9654] = ~(in[375] | in[837]); 
    assign layer_0[9655] = in[805] ^ in[981]; 
    assign layer_0[9656] = in[317] & ~in[477]; 
    assign layer_0[9657] = in[570] & in[667]; 
    assign layer_0[9658] = ~(in[638] ^ in[68]); 
    assign layer_0[9659] = ~in[664] | (in[857] & in[664]); 
    assign layer_0[9660] = ~(in[747] ^ in[221]); 
    assign layer_0[9661] = in[422] ^ in[820]; 
    assign layer_0[9662] = in[34] & ~in[854]; 
    assign layer_0[9663] = ~(in[146] ^ in[468]); 
    assign layer_0[9664] = ~(in[714] ^ in[301]); 
    assign layer_0[9665] = ~in[585] | (in[585] & in[808]); 
    assign layer_0[9666] = ~(in[309] | in[546]); 
    assign layer_0[9667] = in[47]; 
    assign layer_0[9668] = in[730] ^ in[906]; 
    assign layer_0[9669] = in[738] ^ in[177]; 
    assign layer_0[9670] = ~in[993]; 
    assign layer_0[9671] = in[395]; 
    assign layer_0[9672] = ~(in[687] ^ in[362]); 
    assign layer_0[9673] = ~(in[235] & in[969]); 
    assign layer_0[9674] = ~(in[616] & in[968]); 
    assign layer_0[9675] = ~(in[8] & in[177]); 
    assign layer_0[9676] = ~in[441]; 
    assign layer_0[9677] = ~(in[353] ^ in[894]); 
    assign layer_0[9678] = in[811] ^ in[740]; 
    assign layer_0[9679] = in[629]; 
    assign layer_0[9680] = in[225] ^ in[4]; 
    assign layer_0[9681] = ~(in[599] | in[998]); 
    assign layer_0[9682] = ~(in[822] ^ in[662]); 
    assign layer_0[9683] = in[758] ^ in[307]; 
    assign layer_0[9684] = ~(in[300] & in[396]); 
    assign layer_0[9685] = ~(in[325] & in[695]); 
    assign layer_0[9686] = ~in[701] | (in[701] & in[557]); 
    assign layer_0[9687] = ~(in[661] ^ in[663]); 
    assign layer_0[9688] = ~in[245] | (in[350] & in[245]); 
    assign layer_0[9689] = 1'b0; 
    assign layer_0[9690] = ~in[780] | (in[382] & in[780]); 
    assign layer_0[9691] = ~(in[581] & in[969]); 
    assign layer_0[9692] = in[836] ^ in[741]; 
    assign layer_0[9693] = in[498] ^ in[463]; 
    assign layer_0[9694] = in[913] ^ in[131]; 
    assign layer_0[9695] = in[792] | in[580]; 
    assign layer_0[9696] = in[759]; 
    assign layer_0[9697] = in[619] & ~in[825]; 
    assign layer_0[9698] = ~(in[94] ^ in[926]); 
    assign layer_0[9699] = ~(in[690] ^ in[850]); 
    assign layer_0[9700] = ~(in[34] ^ in[877]); 
    assign layer_0[9701] = ~in[297]; 
    assign layer_0[9702] = ~(in[719] | in[589]); 
    assign layer_0[9703] = ~(in[142] ^ in[945]); 
    assign layer_0[9704] = ~(in[614] & in[823]); 
    assign layer_0[9705] = ~(in[766] ^ in[509]); 
    assign layer_0[9706] = ~in[328] | (in[328] & in[398]); 
    assign layer_0[9707] = in[573] ^ in[525]; 
    assign layer_0[9708] = in[661] ^ in[503]; 
    assign layer_0[9709] = in[902] ^ in[942]; 
    assign layer_0[9710] = ~(in[587] | in[924]); 
    assign layer_0[9711] = ~in[588]; 
    assign layer_0[9712] = ~in[267]; 
    assign layer_0[9713] = in[583] ^ in[589]; 
    assign layer_0[9714] = ~(in[478] | in[370]); 
    assign layer_0[9715] = in[539] & ~in[69]; 
    assign layer_0[9716] = in[204] & ~in[781]; 
    assign layer_0[9717] = in[744]; 
    assign layer_0[9718] = in[878] & ~in[512]; 
    assign layer_0[9719] = ~in[501] | (in[501] & in[814]); 
    assign layer_0[9720] = ~in[390] | (in[984] & in[390]); 
    assign layer_0[9721] = in[129] ^ in[788]; 
    assign layer_0[9722] = ~(in[597] ^ in[816]); 
    assign layer_0[9723] = ~in[652]; 
    assign layer_0[9724] = ~(in[619] & in[792]); 
    assign layer_0[9725] = ~(in[241] | in[923]); 
    assign layer_0[9726] = ~(in[989] | in[760]); 
    assign layer_0[9727] = ~in[216] | (in[769] & in[216]); 
    assign layer_0[9728] = ~(in[2] ^ in[536]); 
    assign layer_0[9729] = ~in[634] | (in[634] & in[529]); 
    assign layer_0[9730] = in[160] & ~in[889]; 
    assign layer_0[9731] = ~(in[810] ^ in[858]); 
    assign layer_0[9732] = in[71] & ~in[223]; 
    assign layer_0[9733] = in[372]; 
    assign layer_0[9734] = in[134]; 
    assign layer_0[9735] = in[334] ^ in[537]; 
    assign layer_0[9736] = in[605] ^ in[493]; 
    assign layer_0[9737] = ~in[147] | (in[147] & in[245]); 
    assign layer_0[9738] = ~in[716] | (in[716] & in[875]); 
    assign layer_0[9739] = in[282]; 
    assign layer_0[9740] = in[239]; 
    assign layer_0[9741] = in[711]; 
    assign layer_0[9742] = ~in[228]; 
    assign layer_0[9743] = ~(in[724] ^ in[644]); 
    assign layer_0[9744] = in[506] & ~in[73]; 
    assign layer_0[9745] = ~in[437]; 
    assign layer_0[9746] = in[739]; 
    assign layer_0[9747] = ~(in[520] | in[115]); 
    assign layer_0[9748] = in[915] | in[241]; 
    assign layer_0[9749] = ~(in[329] & in[700]); 
    assign layer_0[9750] = in[904]; 
    assign layer_0[9751] = ~in[194] | (in[194] & in[965]); 
    assign layer_0[9752] = in[983] ^ in[601]; 
    assign layer_0[9753] = ~(in[330] ^ in[647]); 
    assign layer_0[9754] = ~(in[555] ^ in[548]); 
    assign layer_0[9755] = in[380] & in[622]; 
    assign layer_0[9756] = in[550] | in[903]; 
    assign layer_0[9757] = in[602] ^ in[588]; 
    assign layer_0[9758] = in[74] ^ in[708]; 
    assign layer_0[9759] = in[841] | in[512]; 
    assign layer_0[9760] = ~(in[650] ^ in[699]); 
    assign layer_0[9761] = ~(in[958] & in[589]); 
    assign layer_0[9762] = in[265] | in[232]; 
    assign layer_0[9763] = in[238]; 
    assign layer_0[9764] = in[853] ^ in[265]; 
    assign layer_0[9765] = in[412] ^ in[918]; 
    assign layer_0[9766] = ~(in[552] | in[496]); 
    assign layer_0[9767] = in[385] ^ in[596]; 
    assign layer_0[9768] = in[663] & ~in[336]; 
    assign layer_0[9769] = ~in[715]; 
    assign layer_0[9770] = in[441]; 
    assign layer_0[9771] = ~in[679] | (in[679] & in[758]); 
    assign layer_0[9772] = ~in[268] | (in[268] & in[853]); 
    assign layer_0[9773] = ~(in[887] ^ in[886]); 
    assign layer_0[9774] = in[229] & in[399]; 
    assign layer_0[9775] = in[442] & ~in[907]; 
    assign layer_0[9776] = ~(in[144] ^ in[1018]); 
    assign layer_0[9777] = ~(in[733] | in[355]); 
    assign layer_0[9778] = in[63]; 
    assign layer_0[9779] = ~(in[518] & in[377]); 
    assign layer_0[9780] = in[909] & ~in[294]; 
    assign layer_0[9781] = in[965]; 
    assign layer_0[9782] = ~(in[857] ^ in[612]); 
    assign layer_0[9783] = in[275] ^ in[263]; 
    assign layer_0[9784] = in[25]; 
    assign layer_0[9785] = ~in[1003] | (in[659] & in[1003]); 
    assign layer_0[9786] = in[692]; 
    assign layer_0[9787] = ~in[849]; 
    assign layer_0[9788] = ~in[206] | (in[564] & in[206]); 
    assign layer_0[9789] = ~(in[840] ^ in[875]); 
    assign layer_0[9790] = ~in[296]; 
    assign layer_0[9791] = in[632] & ~in[878]; 
    assign layer_0[9792] = ~in[501] | (in[501] & in[731]); 
    assign layer_0[9793] = in[633]; 
    assign layer_0[9794] = ~in[264] | (in[517] & in[264]); 
    assign layer_0[9795] = in[856]; 
    assign layer_0[9796] = in[708] & in[127]; 
    assign layer_0[9797] = ~in[619] | (in[741] & in[619]); 
    assign layer_0[9798] = ~in[706]; 
    assign layer_0[9799] = ~(in[301] ^ in[812]); 
    assign layer_0[9800] = ~(in[838] ^ in[628]); 
    assign layer_0[9801] = ~(in[584] ^ in[458]); 
    assign layer_0[9802] = in[320] & in[642]; 
    assign layer_0[9803] = ~(in[621] ^ in[177]); 
    assign layer_0[9804] = in[210] & ~in[888]; 
    assign layer_0[9805] = ~in[313]; 
    assign layer_0[9806] = ~(in[491] & in[645]); 
    assign layer_0[9807] = ~(in[966] | in[899]); 
    assign layer_0[9808] = ~(in[804] ^ in[924]); 
    assign layer_0[9809] = ~in[627] | (in[887] & in[627]); 
    assign layer_0[9810] = ~in[388] | (in[544] & in[388]); 
    assign layer_0[9811] = in[580] ^ in[179]; 
    assign layer_0[9812] = in[931] | in[326]; 
    assign layer_0[9813] = in[301]; 
    assign layer_0[9814] = in[196] ^ in[4]; 
    assign layer_0[9815] = ~in[340] | (in[340] & in[735]); 
    assign layer_0[9816] = ~(in[910] ^ in[467]); 
    assign layer_0[9817] = ~in[306]; 
    assign layer_0[9818] = in[268]; 
    assign layer_0[9819] = in[885] ^ in[581]; 
    assign layer_0[9820] = in[304]; 
    assign layer_0[9821] = ~in[911]; 
    assign layer_0[9822] = ~(in[263] ^ in[889]); 
    assign layer_0[9823] = ~in[997]; 
    assign layer_0[9824] = in[301] ^ in[316]; 
    assign layer_0[9825] = in[19] & ~in[237]; 
    assign layer_0[9826] = ~(in[80] ^ in[388]); 
    assign layer_0[9827] = in[793] ^ in[997]; 
    assign layer_0[9828] = in[612]; 
    assign layer_0[9829] = ~in[388]; 
    assign layer_0[9830] = ~in[399]; 
    assign layer_0[9831] = in[806]; 
    assign layer_0[9832] = ~in[809]; 
    assign layer_0[9833] = ~(in[906] | in[210]); 
    assign layer_0[9834] = in[956] & ~in[42]; 
    assign layer_0[9835] = in[806] & ~in[702]; 
    assign layer_0[9836] = in[703] & in[833]; 
    assign layer_0[9837] = in[760] & ~in[418]; 
    assign layer_0[9838] = in[49] ^ in[998]; 
    assign layer_0[9839] = in[553] & in[391]; 
    assign layer_0[9840] = in[130] & ~in[585]; 
    assign layer_0[9841] = in[514] | in[324]; 
    assign layer_0[9842] = ~(in[371] | in[937]); 
    assign layer_0[9843] = ~in[236]; 
    assign layer_0[9844] = ~(in[272] & in[881]); 
    assign layer_0[9845] = ~(in[28] & in[551]); 
    assign layer_0[9846] = in[86]; 
    assign layer_0[9847] = ~(in[236] & in[428]); 
    assign layer_0[9848] = in[936] ^ in[616]; 
    assign layer_0[9849] = in[313]; 
    assign layer_0[9850] = ~in[918] | (in[952] & in[918]); 
    assign layer_0[9851] = ~(in[323] | in[562]); 
    assign layer_0[9852] = ~(in[612] ^ in[444]); 
    assign layer_0[9853] = in[839]; 
    assign layer_0[9854] = ~in[925] | (in[925] & in[833]); 
    assign layer_0[9855] = ~(in[749] ^ in[748]); 
    assign layer_0[9856] = in[421] & in[199]; 
    assign layer_0[9857] = in[854] ^ in[704]; 
    assign layer_0[9858] = ~(in[501] | in[260]); 
    assign layer_0[9859] = in[72]; 
    assign layer_0[9860] = in[549] & ~in[674]; 
    assign layer_0[9861] = ~(in[505] | in[976]); 
    assign layer_0[9862] = in[596] & ~in[810]; 
    assign layer_0[9863] = in[933]; 
    assign layer_0[9864] = in[917] ^ in[565]; 
    assign layer_0[9865] = ~(in[570] ^ in[795]); 
    assign layer_0[9866] = in[466]; 
    assign layer_0[9867] = ~(in[686] ^ in[337]); 
    assign layer_0[9868] = ~(in[691] ^ in[946]); 
    assign layer_0[9869] = in[1004] ^ in[314]; 
    assign layer_0[9870] = ~(in[547] | in[340]); 
    assign layer_0[9871] = ~(in[175] & in[112]); 
    assign layer_0[9872] = ~(in[825] & in[151]); 
    assign layer_0[9873] = ~in[51]; 
    assign layer_0[9874] = 1'b1; 
    assign layer_0[9875] = in[220] & ~in[527]; 
    assign layer_0[9876] = ~in[954] | (in[954] & in[220]); 
    assign layer_0[9877] = in[793]; 
    assign layer_0[9878] = in[638] ^ in[82]; 
    assign layer_0[9879] = ~(in[879] | in[598]); 
    assign layer_0[9880] = ~in[564]; 
    assign layer_0[9881] = in[959] ^ in[613]; 
    assign layer_0[9882] = in[71] & ~in[79]; 
    assign layer_0[9883] = in[99]; 
    assign layer_0[9884] = ~(in[699] ^ in[588]); 
    assign layer_0[9885] = ~in[809]; 
    assign layer_0[9886] = ~(in[570] | in[922]); 
    assign layer_0[9887] = in[728]; 
    assign layer_0[9888] = ~in[905] | (in[905] & in[852]); 
    assign layer_0[9889] = in[602] & ~in[541]; 
    assign layer_0[9890] = in[927] ^ in[285]; 
    assign layer_0[9891] = ~(in[176] | in[560]); 
    assign layer_0[9892] = in[938] | in[161]; 
    assign layer_0[9893] = in[821] & in[822]; 
    assign layer_0[9894] = in[924]; 
    assign layer_0[9895] = in[276] & ~in[461]; 
    assign layer_0[9896] = in[572] | in[63]; 
    assign layer_0[9897] = ~in[539]; 
    assign layer_0[9898] = ~(in[461] ^ in[968]); 
    assign layer_0[9899] = ~in[466] | (in[466] & in[14]); 
    assign layer_0[9900] = in[668] | in[683]; 
    assign layer_0[9901] = ~(in[38] | in[918]); 
    assign layer_0[9902] = ~(in[782] ^ in[462]); 
    assign layer_0[9903] = ~(in[714] | in[940]); 
    assign layer_0[9904] = ~(in[133] ^ in[338]); 
    assign layer_0[9905] = ~in[871]; 
    assign layer_0[9906] = in[791] ^ in[604]; 
    assign layer_0[9907] = ~(in[329] ^ in[432]); 
    assign layer_0[9908] = ~in[915]; 
    assign layer_0[9909] = ~in[459]; 
    assign layer_0[9910] = ~in[283] | (in[718] & in[283]); 
    assign layer_0[9911] = ~(in[683] & in[168]); 
    assign layer_0[9912] = ~in[714]; 
    assign layer_0[9913] = ~(in[344] ^ in[574]); 
    assign layer_0[9914] = in[316] | in[274]; 
    assign layer_0[9915] = ~(in[383] ^ in[42]); 
    assign layer_0[9916] = 1'b1; 
    assign layer_0[9917] = in[875] ^ in[564]; 
    assign layer_0[9918] = ~(in[304] ^ in[67]); 
    assign layer_0[9919] = ~in[661]; 
    assign layer_0[9920] = in[324]; 
    assign layer_0[9921] = in[989] ^ in[685]; 
    assign layer_0[9922] = 1'b1; 
    assign layer_0[9923] = in[883] ^ in[899]; 
    assign layer_0[9924] = ~(in[350] | in[384]); 
    assign layer_0[9925] = in[565] & ~in[258]; 
    assign layer_0[9926] = ~(in[616] ^ in[615]); 
    assign layer_0[9927] = in[192] | in[841]; 
    assign layer_0[9928] = ~in[330] | (in[330] & in[903]); 
    assign layer_0[9929] = in[250] & ~in[902]; 
    assign layer_0[9930] = in[253] & in[795]; 
    assign layer_0[9931] = ~(in[928] & in[343]); 
    assign layer_0[9932] = ~in[888]; 
    assign layer_0[9933] = in[84] & ~in[987]; 
    assign layer_0[9934] = in[45] ^ in[40]; 
    assign layer_0[9935] = in[871] ^ in[291]; 
    assign layer_0[9936] = ~in[741] | (in[741] & in[66]); 
    assign layer_0[9937] = in[1015] & ~in[937]; 
    assign layer_0[9938] = ~in[115] | (in[115] & in[881]); 
    assign layer_0[9939] = ~in[233] | (in[273] & in[233]); 
    assign layer_0[9940] = ~in[116] | (in[116] & in[777]); 
    assign layer_0[9941] = ~(in[283] ^ in[333]); 
    assign layer_0[9942] = in[908] | in[994]; 
    assign layer_0[9943] = ~(in[625] ^ in[612]); 
    assign layer_0[9944] = ~(in[760] & in[937]); 
    assign layer_0[9945] = in[680] & ~in[604]; 
    assign layer_0[9946] = in[452]; 
    assign layer_0[9947] = ~(in[124] ^ in[92]); 
    assign layer_0[9948] = in[333] & ~in[239]; 
    assign layer_0[9949] = ~(in[714] ^ in[699]); 
    assign layer_0[9950] = in[616]; 
    assign layer_0[9951] = in[887]; 
    assign layer_0[9952] = in[963] & in[603]; 
    assign layer_0[9953] = ~in[79]; 
    assign layer_0[9954] = ~in[979]; 
    assign layer_0[9955] = ~in[637]; 
    assign layer_0[9956] = ~in[404] | (in[404] & in[843]); 
    assign layer_0[9957] = in[358] & ~in[903]; 
    assign layer_0[9958] = in[609] ^ in[396]; 
    assign layer_0[9959] = ~in[341]; 
    assign layer_0[9960] = in[808] | in[821]; 
    assign layer_0[9961] = in[51]; 
    assign layer_0[9962] = in[667] | in[518]; 
    assign layer_0[9963] = in[43] ^ in[912]; 
    assign layer_0[9964] = ~in[558]; 
    assign layer_0[9965] = ~(in[267] ^ in[444]); 
    assign layer_0[9966] = ~in[12] | (in[815] & in[12]); 
    assign layer_0[9967] = in[683] ^ in[645]; 
    assign layer_0[9968] = in[624] & ~in[675]; 
    assign layer_0[9969] = in[641] ^ in[299]; 
    assign layer_0[9970] = in[615] & in[657]; 
    assign layer_0[9971] = ~in[515]; 
    assign layer_0[9972] = ~in[792]; 
    assign layer_0[9973] = ~(in[1001] ^ in[243]); 
    assign layer_0[9974] = ~(in[6] ^ in[409]); 
    assign layer_0[9975] = ~(in[27] & in[970]); 
    assign layer_0[9976] = 1'b1; 
    assign layer_0[9977] = in[937] & in[118]; 
    assign layer_0[9978] = ~in[174] | (in[174] & in[85]); 
    assign layer_0[9979] = in[959] & in[290]; 
    assign layer_0[9980] = in[754] ^ in[639]; 
    assign layer_0[9981] = in[949] ^ in[244]; 
    assign layer_0[9982] = ~in[377]; 
    assign layer_0[9983] = ~(in[206] | in[664]); 
    assign layer_0[9984] = ~(in[260] | in[948]); 
    assign layer_0[9985] = ~in[378] | (in[860] & in[378]); 
    assign layer_0[9986] = ~in[325]; 
    assign layer_0[9987] = ~(in[483] ^ in[413]); 
    assign layer_0[9988] = ~(in[514] ^ in[759]); 
    assign layer_0[9989] = ~in[699] | (in[873] & in[699]); 
    assign layer_0[9990] = in[716] & ~in[503]; 
    assign layer_0[9991] = ~(in[648] ^ in[568]); 
    assign layer_0[9992] = ~(in[237] ^ in[747]); 
    assign layer_0[9993] = ~in[137] | (in[137] & in[470]); 
    assign layer_0[9994] = ~in[517]; 
    assign layer_0[9995] = in[174] & ~in[527]; 
    assign layer_0[9996] = in[428] & in[484]; 
    assign layer_0[9997] = ~(in[29] | in[570]); 
    assign layer_0[9998] = ~(in[904] ^ in[997]); 
    assign layer_0[9999] = ~(in[417] ^ in[551]); 
    assign layer_0[10000] = in[521] ^ in[69]; 
    assign layer_0[10001] = ~in[60]; 
    assign layer_0[10002] = in[585] ^ in[616]; 
    assign layer_0[10003] = ~(in[241] & in[555]); 
    assign layer_0[10004] = in[691]; 
    assign layer_0[10005] = in[617] ^ in[83]; 
    assign layer_0[10006] = in[865] & in[641]; 
    assign layer_0[10007] = in[933] | in[211]; 
    assign layer_0[10008] = ~(in[677] ^ in[550]); 
    assign layer_0[10009] = 1'b0; 
    assign layer_0[10010] = ~(in[68] | in[732]); 
    assign layer_0[10011] = ~(in[534] & in[35]); 
    assign layer_0[10012] = ~in[569]; 
    assign layer_0[10013] = in[687] & ~in[876]; 
    assign layer_0[10014] = ~(in[388] & in[940]); 
    assign layer_0[10015] = ~in[956]; 
    assign layer_0[10016] = ~(in[54] & in[133]); 
    assign layer_0[10017] = ~(in[38] & in[103]); 
    assign layer_0[10018] = in[449] & in[361]; 
    assign layer_0[10019] = in[377] & in[881]; 
    assign layer_0[10020] = ~(in[17] ^ in[375]); 
    assign layer_0[10021] = ~(in[688] & in[79]); 
    assign layer_0[10022] = ~(in[977] | in[75]); 
    assign layer_0[10023] = in[239] & ~in[366]; 
    assign layer_0[10024] = ~in[175] | (in[175] & in[897]); 
    assign layer_0[10025] = ~in[669]; 
    assign layer_0[10026] = in[75] & ~in[886]; 
    assign layer_0[10027] = in[970]; 
    assign layer_0[10028] = ~in[178] | (in[472] & in[178]); 
    assign layer_0[10029] = in[595] ^ in[355]; 
    assign layer_0[10030] = ~in[997] | (in[997] & in[999]); 
    assign layer_0[10031] = in[450] ^ in[892]; 
    assign layer_0[10032] = ~(in[933] ^ in[324]); 
    assign layer_0[10033] = in[33]; 
    assign layer_0[10034] = ~in[940] | (in[2] & in[940]); 
    assign layer_0[10035] = ~(in[552] ^ in[644]); 
    assign layer_0[10036] = ~(in[395] | in[959]); 
    assign layer_0[10037] = in[604] ^ in[607]; 
    assign layer_0[10038] = in[323] & in[244]; 
    assign layer_0[10039] = in[924] & ~in[504]; 
    assign layer_0[10040] = ~in[471]; 
    assign layer_0[10041] = in[580] & ~in[499]; 
    assign layer_0[10042] = ~in[595]; 
    assign layer_0[10043] = in[650]; 
    assign layer_0[10044] = in[803] | in[193]; 
    assign layer_0[10045] = ~(in[76] & in[786]); 
    assign layer_0[10046] = ~(in[996] ^ in[985]); 
    assign layer_0[10047] = in[115]; 
    assign layer_0[10048] = in[827] | in[904]; 
    assign layer_0[10049] = in[320] & ~in[830]; 
    assign layer_0[10050] = ~in[634] | (in[634] & in[521]); 
    assign layer_0[10051] = in[836] & ~in[745]; 
    assign layer_0[10052] = in[827] & in[9]; 
    assign layer_0[10053] = in[177] | in[895]; 
    assign layer_0[10054] = ~in[892]; 
    assign layer_0[10055] = in[934] & in[827]; 
    assign layer_0[10056] = ~in[651] | (in[883] & in[651]); 
    assign layer_0[10057] = in[994] | in[541]; 
    assign layer_0[10058] = ~(in[776] ^ in[1015]); 
    assign layer_0[10059] = in[291]; 
    assign layer_0[10060] = in[142]; 
    assign layer_0[10061] = ~in[76] | (in[76] & in[673]); 
    assign layer_0[10062] = ~in[83]; 
    assign layer_0[10063] = ~in[747]; 
    assign layer_0[10064] = ~(in[200] & in[889]); 
    assign layer_0[10065] = in[311] ^ in[656]; 
    assign layer_0[10066] = in[537] & in[437]; 
    assign layer_0[10067] = ~(in[227] ^ in[642]); 
    assign layer_0[10068] = ~(in[983] ^ in[985]); 
    assign layer_0[10069] = ~(in[695] ^ in[919]); 
    assign layer_0[10070] = ~(in[744] & in[611]); 
    assign layer_0[10071] = in[429]; 
    assign layer_0[10072] = ~(in[897] ^ in[585]); 
    assign layer_0[10073] = in[796] & ~in[907]; 
    assign layer_0[10074] = ~in[525] | (in[525] & in[949]); 
    assign layer_0[10075] = in[589] ^ in[402]; 
    assign layer_0[10076] = in[408] & in[8]; 
    assign layer_0[10077] = ~in[412]; 
    assign layer_0[10078] = in[486] ^ in[845]; 
    assign layer_0[10079] = ~(in[64] | in[1022]); 
    assign layer_0[10080] = in[83] & in[301]; 
    assign layer_0[10081] = in[757] ^ in[312]; 
    assign layer_0[10082] = in[881] ^ in[22]; 
    assign layer_0[10083] = ~(in[619] ^ in[499]); 
    assign layer_0[10084] = in[387] & ~in[351]; 
    assign layer_0[10085] = ~in[934]; 
    assign layer_0[10086] = in[326] ^ in[602]; 
    assign layer_0[10087] = in[917] ^ in[434]; 
    assign layer_0[10088] = ~in[782] | (in[151] & in[782]); 
    assign layer_0[10089] = in[650] & ~in[807]; 
    assign layer_0[10090] = ~in[35] | (in[1005] & in[35]); 
    assign layer_0[10091] = ~in[1010]; 
    assign layer_0[10092] = in[307] & ~in[788]; 
    assign layer_0[10093] = in[812] & ~in[1007]; 
    assign layer_0[10094] = ~(in[930] ^ in[735]); 
    assign layer_0[10095] = in[538] ^ in[585]; 
    assign layer_0[10096] = in[955] ^ in[739]; 
    assign layer_0[10097] = in[678]; 
    assign layer_0[10098] = in[1010] | in[981]; 
    assign layer_0[10099] = ~(in[808] ^ in[809]); 
    assign layer_0[10100] = ~in[281]; 
    assign layer_0[10101] = ~(in[283] | in[285]); 
    assign layer_0[10102] = in[312] & ~in[639]; 
    assign layer_0[10103] = in[262] ^ in[469]; 
    assign layer_0[10104] = ~in[795]; 
    assign layer_0[10105] = in[635] & ~in[219]; 
    assign layer_0[10106] = ~(in[412] | in[718]); 
    assign layer_0[10107] = in[893]; 
    assign layer_0[10108] = in[354] ^ in[841]; 
    assign layer_0[10109] = 1'b0; 
    assign layer_0[10110] = ~(in[109] ^ in[538]); 
    assign layer_0[10111] = in[276] & ~in[673]; 
    assign layer_0[10112] = in[427]; 
    assign layer_0[10113] = 1'b0; 
    assign layer_0[10114] = ~in[517] | (in[517] & in[611]); 
    assign layer_0[10115] = in[963] ^ in[597]; 
    assign layer_0[10116] = ~(in[954] | in[206]); 
    assign layer_0[10117] = in[465]; 
    assign layer_0[10118] = in[638] ^ in[610]; 
    assign layer_0[10119] = in[28]; 
    assign layer_0[10120] = in[404]; 
    assign layer_0[10121] = ~(in[811] | in[46]); 
    assign layer_0[10122] = in[12] ^ in[792]; 
    assign layer_0[10123] = ~in[388]; 
    assign layer_0[10124] = ~in[29]; 
    assign layer_0[10125] = ~(in[437] ^ in[379]); 
    assign layer_0[10126] = ~in[663] | (in[663] & in[502]); 
    assign layer_0[10127] = ~(in[338] ^ in[501]); 
    assign layer_0[10128] = in[953] ^ in[603]; 
    assign layer_0[10129] = ~in[700] | (in[304] & in[700]); 
    assign layer_0[10130] = in[997] | in[321]; 
    assign layer_0[10131] = ~(in[353] ^ in[608]); 
    assign layer_0[10132] = in[454]; 
    assign layer_0[10133] = ~in[167] | (in[592] & in[167]); 
    assign layer_0[10134] = ~(in[807] ^ in[350]); 
    assign layer_0[10135] = in[953] ^ in[226]; 
    assign layer_0[10136] = ~(in[427] ^ in[301]); 
    assign layer_0[10137] = in[651] ^ in[876]; 
    assign layer_0[10138] = ~in[109] | (in[109] & in[488]); 
    assign layer_0[10139] = in[942]; 
    assign layer_0[10140] = ~(in[889] ^ in[950]); 
    assign layer_0[10141] = ~in[948]; 
    assign layer_0[10142] = ~(in[878] ^ in[698]); 
    assign layer_0[10143] = 1'b0; 
    assign layer_0[10144] = ~in[887]; 
    assign layer_0[10145] = ~in[618]; 
    assign layer_0[10146] = ~in[469] | (in[469] & in[643]); 
    assign layer_0[10147] = in[793] | in[811]; 
    assign layer_0[10148] = ~(in[715] & in[484]); 
    assign layer_0[10149] = in[371] & ~in[503]; 
    assign layer_0[10150] = ~in[309]; 
    assign layer_0[10151] = ~(in[482] | in[606]); 
    assign layer_0[10152] = ~in[424] | (in[268] & in[424]); 
    assign layer_0[10153] = in[744] ^ in[955]; 
    assign layer_0[10154] = ~(in[844] & in[323]); 
    assign layer_0[10155] = in[904] & ~in[80]; 
    assign layer_0[10156] = in[759]; 
    assign layer_0[10157] = in[825]; 
    assign layer_0[10158] = in[673] | in[29]; 
    assign layer_0[10159] = in[97] ^ in[884]; 
    assign layer_0[10160] = in[1000] | in[289]; 
    assign layer_0[10161] = in[202] ^ in[101]; 
    assign layer_0[10162] = in[620] ^ in[279]; 
    assign layer_0[10163] = ~(in[842] | in[837]); 
    assign layer_0[10164] = in[635] & in[650]; 
    assign layer_0[10165] = ~in[872]; 
    assign layer_0[10166] = ~in[334]; 
    assign layer_0[10167] = ~in[997] | (in[517] & in[997]); 
    assign layer_0[10168] = ~(in[963] ^ in[195]); 
    assign layer_0[10169] = ~(in[1016] & in[985]); 
    assign layer_0[10170] = in[937] ^ in[757]; 
    assign layer_0[10171] = in[332] ^ in[124]; 
    assign layer_0[10172] = in[420] & ~in[584]; 
    assign layer_0[10173] = in[177] ^ in[507]; 
    assign layer_0[10174] = ~(in[365] ^ in[49]); 
    assign layer_0[10175] = in[598] | in[302]; 
    assign layer_0[10176] = ~(in[289] | in[829]); 
    assign layer_0[10177] = ~in[539]; 
    assign layer_0[10178] = in[249] & ~in[470]; 
    assign layer_0[10179] = ~in[920] | (in[964] & in[920]); 
    assign layer_0[10180] = in[493] ^ in[283]; 
    assign layer_0[10181] = ~(in[533] ^ in[870]); 
    assign layer_0[10182] = ~(in[590] & in[906]); 
    assign layer_0[10183] = ~(in[100] ^ in[148]); 
    assign layer_0[10184] = in[566] | in[565]; 
    assign layer_0[10185] = ~(in[588] | in[729]); 
    assign layer_0[10186] = in[461]; 
    assign layer_0[10187] = ~in[821]; 
    assign layer_0[10188] = ~in[63]; 
    assign layer_0[10189] = in[218] | in[656]; 
    assign layer_0[10190] = in[934] ^ in[698]; 
    assign layer_0[10191] = in[173] ^ in[819]; 
    assign layer_0[10192] = in[961] ^ in[1002]; 
    assign layer_0[10193] = ~(in[214] & in[616]); 
    assign layer_0[10194] = ~(in[294] ^ in[462]); 
    assign layer_0[10195] = in[175] & ~in[322]; 
    assign layer_0[10196] = ~(in[295] & in[122]); 
    assign layer_0[10197] = in[651] & ~in[229]; 
    assign layer_0[10198] = in[612] ^ in[581]; 
    assign layer_0[10199] = ~(in[353] ^ in[481]); 
    assign layer_0[10200] = ~in[276] | (in[755] & in[276]); 
    assign layer_0[10201] = in[1002]; 
    assign layer_0[10202] = in[744]; 
    assign layer_0[10203] = ~(in[163] ^ in[918]); 
    assign layer_0[10204] = in[760]; 
    assign layer_0[10205] = in[100] & ~in[30]; 
    assign layer_0[10206] = in[539] ^ in[139]; 
    assign layer_0[10207] = ~in[488] | (in[488] & in[854]); 
    assign layer_0[10208] = ~in[842]; 
    assign layer_0[10209] = ~in[481] | (in[481] & in[580]); 
    assign layer_0[10210] = in[837] ^ in[504]; 
    assign layer_0[10211] = in[568] & ~in[903]; 
    assign layer_0[10212] = ~(in[775] | in[336]); 
    assign layer_0[10213] = in[19] & ~in[232]; 
    assign layer_0[10214] = in[633] & ~in[66]; 
    assign layer_0[10215] = ~(in[886] ^ in[349]); 
    assign layer_0[10216] = ~(in[50] ^ in[822]); 
    assign layer_0[10217] = in[891] ^ in[727]; 
    assign layer_0[10218] = in[467] & ~in[891]; 
    assign layer_0[10219] = ~in[137]; 
    assign layer_0[10220] = ~in[518]; 
    assign layer_0[10221] = in[132]; 
    assign layer_0[10222] = in[436]; 
    assign layer_0[10223] = ~in[27] | (in[547] & in[27]); 
    assign layer_0[10224] = in[966] & in[965]; 
    assign layer_0[10225] = ~(in[315] ^ in[477]); 
    assign layer_0[10226] = ~in[8] | (in[8] & in[840]); 
    assign layer_0[10227] = ~in[84] | (in[62] & in[84]); 
    assign layer_0[10228] = ~in[518]; 
    assign layer_0[10229] = ~in[250] | (in[560] & in[250]); 
    assign layer_0[10230] = ~(in[631] ^ in[874]); 
    assign layer_0[10231] = in[518] & ~in[984]; 
    assign layer_0[10232] = ~(in[890] | in[13]); 
    assign layer_0[10233] = ~(in[537] ^ in[520]); 
    assign layer_0[10234] = in[12] ^ in[170]; 
    assign layer_0[10235] = in[552] ^ in[753]; 
    assign layer_0[10236] = in[200] & ~in[574]; 
    assign layer_0[10237] = in[302] & ~in[786]; 
    assign layer_0[10238] = ~(in[470] & in[132]); 
    assign layer_0[10239] = in[725] | in[255]; 
    assign layer_0[10240] = ~(in[537] ^ in[109]); 
    assign layer_0[10241] = in[50]; 
    assign layer_0[10242] = ~(in[812] | in[336]); 
    assign layer_0[10243] = in[706] & ~in[473]; 
    assign layer_0[10244] = in[140] & ~in[620]; 
    assign layer_0[10245] = ~(in[966] ^ in[998]); 
    assign layer_0[10246] = ~in[457] | (in[457] & in[272]); 
    assign layer_0[10247] = in[393] & ~in[764]; 
    assign layer_0[10248] = in[879] ^ in[626]; 
    assign layer_0[10249] = in[649] ^ in[569]; 
    assign layer_0[10250] = in[475]; 
    assign layer_0[10251] = in[69] ^ in[645]; 
    assign layer_0[10252] = in[244] | in[857]; 
    assign layer_0[10253] = ~(in[848] | in[353]); 
    assign layer_0[10254] = ~in[630]; 
    assign layer_0[10255] = in[286] & ~in[487]; 
    assign layer_0[10256] = in[853] ^ in[634]; 
    assign layer_0[10257] = ~(in[352] ^ in[725]); 
    assign layer_0[10258] = in[673] ^ in[381]; 
    assign layer_0[10259] = in[69] & ~in[821]; 
    assign layer_0[10260] = in[842] | in[499]; 
    assign layer_0[10261] = in[899] ^ in[96]; 
    assign layer_0[10262] = in[804] & ~in[914]; 
    assign layer_0[10263] = ~(in[963] ^ in[584]); 
    assign layer_0[10264] = in[490]; 
    assign layer_0[10265] = in[122] & ~in[629]; 
    assign layer_0[10266] = ~in[127]; 
    assign layer_0[10267] = in[217] ^ in[500]; 
    assign layer_0[10268] = ~in[173]; 
    assign layer_0[10269] = in[857] & ~in[948]; 
    assign layer_0[10270] = in[884] & ~in[123]; 
    assign layer_0[10271] = in[231] ^ in[19]; 
    assign layer_0[10272] = ~(in[477] | in[618]); 
    assign layer_0[10273] = ~(in[89] & in[985]); 
    assign layer_0[10274] = ~(in[838] ^ in[997]); 
    assign layer_0[10275] = ~(in[462] & in[988]); 
    assign layer_0[10276] = ~(in[661] ^ in[569]); 
    assign layer_0[10277] = in[855] ^ in[57]; 
    assign layer_0[10278] = ~in[332] | (in[332] & in[534]); 
    assign layer_0[10279] = in[574] | in[261]; 
    assign layer_0[10280] = ~(in[920] ^ in[883]); 
    assign layer_0[10281] = in[372] ^ in[590]; 
    assign layer_0[10282] = 1'b1; 
    assign layer_0[10283] = ~(in[521] ^ in[222]); 
    assign layer_0[10284] = ~(in[71] | in[875]); 
    assign layer_0[10285] = ~in[595]; 
    assign layer_0[10286] = in[807] ^ in[805]; 
    assign layer_0[10287] = ~in[838]; 
    assign layer_0[10288] = in[503] ^ in[501]; 
    assign layer_0[10289] = ~(in[638] & in[179]); 
    assign layer_0[10290] = ~(in[161] ^ in[989]); 
    assign layer_0[10291] = in[330]; 
    assign layer_0[10292] = ~in[552]; 
    assign layer_0[10293] = in[340] & ~in[660]; 
    assign layer_0[10294] = ~in[574] | (in[574] & in[26]); 
    assign layer_0[10295] = in[115] & in[46]; 
    assign layer_0[10296] = in[203]; 
    assign layer_0[10297] = in[255] & in[487]; 
    assign layer_0[10298] = in[113]; 
    assign layer_0[10299] = ~in[173]; 
    assign layer_0[10300] = ~in[42] | (in[644] & in[42]); 
    assign layer_0[10301] = in[598] ^ in[968]; 
    assign layer_0[10302] = in[307] & in[915]; 
    assign layer_0[10303] = in[732]; 
    assign layer_0[10304] = in[62] | in[878]; 
    assign layer_0[10305] = ~(in[934] ^ in[660]); 
    assign layer_0[10306] = ~(in[975] ^ in[11]); 
    assign layer_0[10307] = 1'b0; 
    assign layer_0[10308] = ~(in[35] | in[880]); 
    assign layer_0[10309] = in[534] & in[584]; 
    assign layer_0[10310] = in[177]; 
    assign layer_0[10311] = in[6] & in[949]; 
    assign layer_0[10312] = in[276] ^ in[261]; 
    assign layer_0[10313] = ~in[464]; 
    assign layer_0[10314] = 1'b1; 
    assign layer_0[10315] = in[545]; 
    assign layer_0[10316] = ~in[1004] | (in[1004] & in[209]); 
    assign layer_0[10317] = ~(in[692] ^ in[724]); 
    assign layer_0[10318] = ~(in[856] ^ in[932]); 
    assign layer_0[10319] = in[333] ^ in[324]; 
    assign layer_0[10320] = in[917] ^ in[208]; 
    assign layer_0[10321] = ~in[820] | (in[820] & in[402]); 
    assign layer_0[10322] = in[908] & ~in[49]; 
    assign layer_0[10323] = ~(in[278] ^ in[656]); 
    assign layer_0[10324] = ~in[328] | (in[328] & in[950]); 
    assign layer_0[10325] = in[720] ^ in[926]; 
    assign layer_0[10326] = ~in[48] | (in[48] & in[273]); 
    assign layer_0[10327] = in[739] | in[639]; 
    assign layer_0[10328] = ~in[904] | (in[953] & in[904]); 
    assign layer_0[10329] = ~(in[980] ^ in[338]); 
    assign layer_0[10330] = 1'b0; 
    assign layer_0[10331] = ~(in[535] ^ in[656]); 
    assign layer_0[10332] = ~(in[925] | in[868]); 
    assign layer_0[10333] = ~in[695]; 
    assign layer_0[10334] = ~(in[817] ^ in[715]); 
    assign layer_0[10335] = ~in[589]; 
    assign layer_0[10336] = in[60] & ~in[46]; 
    assign layer_0[10337] = ~in[619] | (in[619] & in[792]); 
    assign layer_0[10338] = ~in[388] | (in[786] & in[388]); 
    assign layer_0[10339] = ~(in[519] ^ in[534]); 
    assign layer_0[10340] = ~in[999]; 
    assign layer_0[10341] = in[261] ^ in[264]; 
    assign layer_0[10342] = ~in[331] | (in[331] & in[744]); 
    assign layer_0[10343] = ~(in[489] ^ in[64]); 
    assign layer_0[10344] = ~(in[877] ^ in[292]); 
    assign layer_0[10345] = in[54]; 
    assign layer_0[10346] = in[531] ^ in[330]; 
    assign layer_0[10347] = in[538] & ~in[520]; 
    assign layer_0[10348] = ~in[63] | (in[63] & in[918]); 
    assign layer_0[10349] = ~(in[242] ^ in[913]); 
    assign layer_0[10350] = in[254] & ~in[829]; 
    assign layer_0[10351] = ~in[19]; 
    assign layer_0[10352] = ~in[754]; 
    assign layer_0[10353] = ~in[273] | (in[297] & in[273]); 
    assign layer_0[10354] = ~in[917]; 
    assign layer_0[10355] = ~in[999] | (in[517] & in[999]); 
    assign layer_0[10356] = ~in[128] | (in[128] & in[448]); 
    assign layer_0[10357] = in[400] ^ in[445]; 
    assign layer_0[10358] = in[193] & ~in[352]; 
    assign layer_0[10359] = in[427] & in[919]; 
    assign layer_0[10360] = ~in[132] | (in[132] & in[740]); 
    assign layer_0[10361] = ~(in[73] ^ in[269]); 
    assign layer_0[10362] = ~in[263] | (in[354] & in[263]); 
    assign layer_0[10363] = ~(in[617] ^ in[804]); 
    assign layer_0[10364] = in[619] ^ in[565]; 
    assign layer_0[10365] = in[86] & ~in[142]; 
    assign layer_0[10366] = ~in[890] | (in[798] & in[890]); 
    assign layer_0[10367] = ~(in[521] ^ in[943]); 
    assign layer_0[10368] = ~(in[739] & in[899]); 
    assign layer_0[10369] = in[1009]; 
    assign layer_0[10370] = ~(in[209] & in[469]); 
    assign layer_0[10371] = ~(in[914] ^ in[950]); 
    assign layer_0[10372] = in[295] & in[265]; 
    assign layer_0[10373] = in[2] | in[893]; 
    assign layer_0[10374] = in[362] ^ in[667]; 
    assign layer_0[10375] = in[146] & ~in[715]; 
    assign layer_0[10376] = in[380] & in[851]; 
    assign layer_0[10377] = ~(in[874] ^ in[630]); 
    assign layer_0[10378] = ~(in[129] | in[711]); 
    assign layer_0[10379] = ~in[796] | (in[796] & in[209]); 
    assign layer_0[10380] = in[610] ^ in[518]; 
    assign layer_0[10381] = in[83]; 
    assign layer_0[10382] = in[900] ^ in[842]; 
    assign layer_0[10383] = ~in[507] | (in[302] & in[507]); 
    assign layer_0[10384] = in[818]; 
    assign layer_0[10385] = ~in[739] | (in[814] & in[739]); 
    assign layer_0[10386] = ~(in[554] ^ in[333]); 
    assign layer_0[10387] = in[677] & ~in[930]; 
    assign layer_0[10388] = ~(in[471] ^ in[860]); 
    assign layer_0[10389] = ~(in[736] | in[78]); 
    assign layer_0[10390] = ~(in[984] ^ in[663]); 
    assign layer_0[10391] = ~(in[266] | in[261]); 
    assign layer_0[10392] = in[538] ^ in[233]; 
    assign layer_0[10393] = ~in[433] | (in[433] & in[789]); 
    assign layer_0[10394] = in[634] ^ in[621]; 
    assign layer_0[10395] = in[655]; 
    assign layer_0[10396] = in[92] ^ in[874]; 
    assign layer_0[10397] = ~in[697]; 
    assign layer_0[10398] = ~in[78] | (in[732] & in[78]); 
    assign layer_0[10399] = ~in[243] | (in[243] & in[33]); 
    assign layer_0[10400] = in[502] ^ in[292]; 
    assign layer_0[10401] = ~in[508] | (in[508] & in[344]); 
    assign layer_0[10402] = ~(in[283] ^ in[648]); 
    assign layer_0[10403] = ~in[197] | (in[197] & in[242]); 
    assign layer_0[10404] = 1'b0; 
    assign layer_0[10405] = in[674] ^ in[717]; 
    assign layer_0[10406] = in[458] & ~in[1002]; 
    assign layer_0[10407] = ~(in[564] & in[744]); 
    assign layer_0[10408] = ~in[29] | (in[29] & in[126]); 
    assign layer_0[10409] = in[664] & ~in[952]; 
    assign layer_0[10410] = in[967] & ~in[539]; 
    assign layer_0[10411] = ~in[916] | (in[916] & in[353]); 
    assign layer_0[10412] = ~(in[452] ^ in[449]); 
    assign layer_0[10413] = ~(in[317] ^ in[520]); 
    assign layer_0[10414] = in[396] & in[632]; 
    assign layer_0[10415] = ~in[619] | (in[619] & in[114]); 
    assign layer_0[10416] = in[486] ^ in[109]; 
    assign layer_0[10417] = in[631] & ~in[764]; 
    assign layer_0[10418] = ~(in[709] ^ in[178]); 
    assign layer_0[10419] = ~(in[847] | in[618]); 
    assign layer_0[10420] = ~in[324]; 
    assign layer_0[10421] = ~(in[942] | in[838]); 
    assign layer_0[10422] = in[252] ^ in[34]; 
    assign layer_0[10423] = ~in[787]; 
    assign layer_0[10424] = ~(in[19] | in[1017]); 
    assign layer_0[10425] = in[275]; 
    assign layer_0[10426] = in[853] & ~in[856]; 
    assign layer_0[10427] = in[903] ^ in[842]; 
    assign layer_0[10428] = ~(in[142] & in[663]); 
    assign layer_0[10429] = in[355] & ~in[725]; 
    assign layer_0[10430] = ~(in[807] ^ in[567]); 
    assign layer_0[10431] = ~(in[523] ^ in[671]); 
    assign layer_0[10432] = in[54] & in[357]; 
    assign layer_0[10433] = ~(in[269] & in[811]); 
    assign layer_0[10434] = in[396] & in[894]; 
    assign layer_0[10435] = ~in[630] | (in[986] & in[630]); 
    assign layer_0[10436] = in[500]; 
    assign layer_0[10437] = ~(in[10] ^ in[94]); 
    assign layer_0[10438] = ~in[756]; 
    assign layer_0[10439] = ~(in[870] ^ in[519]); 
    assign layer_0[10440] = ~in[97] | (in[97] & in[870]); 
    assign layer_0[10441] = in[207] ^ in[114]; 
    assign layer_0[10442] = in[35] & ~in[837]; 
    assign layer_0[10443] = ~(in[755] ^ in[497]); 
    assign layer_0[10444] = in[696] & ~in[1014]; 
    assign layer_0[10445] = ~(in[245] ^ in[793]); 
    assign layer_0[10446] = in[944] & in[458]; 
    assign layer_0[10447] = in[211]; 
    assign layer_0[10448] = in[901]; 
    assign layer_0[10449] = ~in[714] | (in[661] & in[714]); 
    assign layer_0[10450] = in[722] & ~in[896]; 
    assign layer_0[10451] = ~(in[878] | in[792]); 
    assign layer_0[10452] = ~in[854] | (in[854] & in[662]); 
    assign layer_0[10453] = in[251]; 
    assign layer_0[10454] = ~in[952] | (in[952] & in[865]); 
    assign layer_0[10455] = ~(in[597] & in[565]); 
    assign layer_0[10456] = in[662]; 
    assign layer_0[10457] = in[225] | in[307]; 
    assign layer_0[10458] = ~(in[687] & in[877]); 
    assign layer_0[10459] = ~(in[292] | in[604]); 
    assign layer_0[10460] = in[134] & ~in[723]; 
    assign layer_0[10461] = in[891] & ~in[829]; 
    assign layer_0[10462] = in[206] ^ in[349]; 
    assign layer_0[10463] = in[446] & in[410]; 
    assign layer_0[10464] = ~(in[294] ^ in[580]); 
    assign layer_0[10465] = ~in[79] | (in[79] & in[917]); 
    assign layer_0[10466] = in[922] & in[717]; 
    assign layer_0[10467] = ~(in[571] ^ in[580]); 
    assign layer_0[10468] = in[702] & ~in[266]; 
    assign layer_0[10469] = in[912] ^ in[419]; 
    assign layer_0[10470] = in[889] ^ in[958]; 
    assign layer_0[10471] = ~(in[467] ^ in[21]); 
    assign layer_0[10472] = in[506] ^ in[982]; 
    assign layer_0[10473] = ~(in[95] ^ in[316]); 
    assign layer_0[10474] = in[136] & ~in[838]; 
    assign layer_0[10475] = in[493] & ~in[816]; 
    assign layer_0[10476] = ~(in[604] & in[84]); 
    assign layer_0[10477] = ~(in[174] ^ in[825]); 
    assign layer_0[10478] = ~in[399]; 
    assign layer_0[10479] = ~(in[408] | in[80]); 
    assign layer_0[10480] = in[557] & ~in[392]; 
    assign layer_0[10481] = ~(in[35] | in[889]); 
    assign layer_0[10482] = ~(in[671] ^ in[74]); 
    assign layer_0[10483] = in[550] ^ in[998]; 
    assign layer_0[10484] = ~(in[760] ^ in[372]); 
    assign layer_0[10485] = in[172] ^ in[326]; 
    assign layer_0[10486] = in[650] ^ in[175]; 
    assign layer_0[10487] = in[507] & ~in[936]; 
    assign layer_0[10488] = in[581] & ~in[790]; 
    assign layer_0[10489] = in[4] & in[267]; 
    assign layer_0[10490] = in[427]; 
    assign layer_0[10491] = ~(in[859] & in[549]); 
    assign layer_0[10492] = in[120] & ~in[507]; 
    assign layer_0[10493] = in[980] ^ in[586]; 
    assign layer_0[10494] = ~in[824]; 
    assign layer_0[10495] = ~(in[554] ^ in[781]); 
    assign layer_0[10496] = in[688] ^ in[911]; 
    assign layer_0[10497] = in[533] | in[309]; 
    assign layer_0[10498] = in[678] ^ in[33]; 
    assign layer_0[10499] = in[909] & in[466]; 
    assign layer_0[10500] = in[949] ^ in[725]; 
    assign layer_0[10501] = ~in[51]; 
    assign layer_0[10502] = ~(in[983] | in[985]); 
    assign layer_0[10503] = ~in[100] | (in[942] & in[100]); 
    assign layer_0[10504] = ~(in[553] ^ in[582]); 
    assign layer_0[10505] = ~in[843] | (in[843] & in[39]); 
    assign layer_0[10506] = in[659] & ~in[657]; 
    assign layer_0[10507] = ~(in[609] ^ in[488]); 
    assign layer_0[10508] = ~(in[902] ^ in[904]); 
    assign layer_0[10509] = ~in[664] | (in[515] & in[664]); 
    assign layer_0[10510] = in[916] ^ in[211]; 
    assign layer_0[10511] = ~(in[715] ^ in[760]); 
    assign layer_0[10512] = in[554] ^ in[918]; 
    assign layer_0[10513] = in[715] & ~in[684]; 
    assign layer_0[10514] = in[786] & ~in[784]; 
    assign layer_0[10515] = ~in[810] | (in[520] & in[810]); 
    assign layer_0[10516] = in[932] ^ in[575]; 
    assign layer_0[10517] = ~in[975] | (in[18] & in[975]); 
    assign layer_0[10518] = in[43] ^ in[669]; 
    assign layer_0[10519] = ~(in[45] ^ in[603]); 
    assign layer_0[10520] = in[310] ^ in[896]; 
    assign layer_0[10521] = in[776] & ~in[260]; 
    assign layer_0[10522] = ~(in[292] ^ in[507]); 
    assign layer_0[10523] = ~(in[47] & in[652]); 
    assign layer_0[10524] = in[930] ^ in[824]; 
    assign layer_0[10525] = in[528]; 
    assign layer_0[10526] = ~(in[549] ^ in[997]); 
    assign layer_0[10527] = ~(in[846] | in[623]); 
    assign layer_0[10528] = in[709] ^ in[732]; 
    assign layer_0[10529] = ~(in[99] | in[540]); 
    assign layer_0[10530] = in[566] ^ in[923]; 
    assign layer_0[10531] = ~(in[761] ^ in[218]); 
    assign layer_0[10532] = ~(in[377] ^ in[728]); 
    assign layer_0[10533] = in[536] ^ in[614]; 
    assign layer_0[10534] = in[476] ^ in[869]; 
    assign layer_0[10535] = ~in[164] | (in[63] & in[164]); 
    assign layer_0[10536] = ~(in[177] ^ in[805]); 
    assign layer_0[10537] = in[451] & ~in[144]; 
    assign layer_0[10538] = in[76] & ~in[810]; 
    assign layer_0[10539] = in[587] & in[231]; 
    assign layer_0[10540] = in[909]; 
    assign layer_0[10541] = in[155] & ~in[759]; 
    assign layer_0[10542] = ~in[118] | (in[788] & in[118]); 
    assign layer_0[10543] = in[452] & in[812]; 
    assign layer_0[10544] = in[876] & ~in[610]; 
    assign layer_0[10545] = ~in[97]; 
    assign layer_0[10546] = in[169] | in[906]; 
    assign layer_0[10547] = in[265] & ~in[885]; 
    assign layer_0[10548] = ~(in[9] ^ in[284]); 
    assign layer_0[10549] = in[404] ^ in[792]; 
    assign layer_0[10550] = ~(in[5] ^ in[884]); 
    assign layer_0[10551] = in[818] | in[1000]; 
    assign layer_0[10552] = ~(in[938] | in[383]); 
    assign layer_0[10553] = ~(in[971] ^ in[651]); 
    assign layer_0[10554] = ~(in[628] & in[910]); 
    assign layer_0[10555] = ~(in[832] | in[486]); 
    assign layer_0[10556] = ~in[935] | (in[953] & in[935]); 
    assign layer_0[10557] = ~(in[694] & in[811]); 
    assign layer_0[10558] = ~(in[451] ^ in[603]); 
    assign layer_0[10559] = ~(in[837] | in[533]); 
    assign layer_0[10560] = in[950] ^ in[919]; 
    assign layer_0[10561] = in[155] & ~in[873]; 
    assign layer_0[10562] = ~(in[466] & in[11]); 
    assign layer_0[10563] = in[4]; 
    assign layer_0[10564] = ~(in[507] & in[759]); 
    assign layer_0[10565] = in[1002] & ~in[693]; 
    assign layer_0[10566] = ~(in[928] | in[739]); 
    assign layer_0[10567] = ~(in[723] & in[920]); 
    assign layer_0[10568] = ~in[121]; 
    assign layer_0[10569] = in[485] & in[89]; 
    assign layer_0[10570] = ~(in[434] ^ in[202]); 
    assign layer_0[10571] = ~(in[381] ^ in[442]); 
    assign layer_0[10572] = in[841]; 
    assign layer_0[10573] = ~in[373] | (in[763] & in[373]); 
    assign layer_0[10574] = ~in[96]; 
    assign layer_0[10575] = in[985] ^ in[764]; 
    assign layer_0[10576] = in[705] & ~in[981]; 
    assign layer_0[10577] = in[290] & in[477]; 
    assign layer_0[10578] = ~(in[587] ^ in[927]); 
    assign layer_0[10579] = in[823] & ~in[820]; 
    assign layer_0[10580] = in[601]; 
    assign layer_0[10581] = ~in[348] | (in[858] & in[348]); 
    assign layer_0[10582] = ~in[788]; 
    assign layer_0[10583] = ~in[850]; 
    assign layer_0[10584] = ~(in[594] ^ in[348]); 
    assign layer_0[10585] = ~(in[694] ^ in[585]); 
    assign layer_0[10586] = ~in[937]; 
    assign layer_0[10587] = in[62] ^ in[461]; 
    assign layer_0[10588] = ~(in[828] | in[547]); 
    assign layer_0[10589] = in[483] ^ in[205]; 
    assign layer_0[10590] = in[879] & in[931]; 
    assign layer_0[10591] = in[532] ^ in[870]; 
    assign layer_0[10592] = in[948]; 
    assign layer_0[10593] = ~(in[957] | in[725]); 
    assign layer_0[10594] = ~(in[995] ^ in[88]); 
    assign layer_0[10595] = in[689] ^ in[808]; 
    assign layer_0[10596] = in[150]; 
    assign layer_0[10597] = ~(in[885] ^ in[909]); 
    assign layer_0[10598] = ~(in[158] & in[860]); 
    assign layer_0[10599] = ~in[936] | (in[977] & in[936]); 
    assign layer_0[10600] = in[188]; 
    assign layer_0[10601] = ~in[830] | (in[830] & in[284]); 
    assign layer_0[10602] = in[908]; 
    assign layer_0[10603] = ~in[389] | (in[389] & in[60]); 
    assign layer_0[10604] = ~(in[999] | in[749]); 
    assign layer_0[10605] = in[652] & ~in[76]; 
    assign layer_0[10606] = in[604] ^ in[600]; 
    assign layer_0[10607] = in[622] ^ in[730]; 
    assign layer_0[10608] = in[518]; 
    assign layer_0[10609] = in[932] ^ in[461]; 
    assign layer_0[10610] = 1'b1; 
    assign layer_0[10611] = in[105]; 
    assign layer_0[10612] = in[726] & ~in[51]; 
    assign layer_0[10613] = in[175] | in[127]; 
    assign layer_0[10614] = in[263] & in[326]; 
    assign layer_0[10615] = in[764] & ~in[636]; 
    assign layer_0[10616] = in[929] ^ in[924]; 
    assign layer_0[10617] = ~in[463]; 
    assign layer_0[10618] = ~(in[872] ^ in[598]); 
    assign layer_0[10619] = ~(in[904] ^ in[876]); 
    assign layer_0[10620] = ~in[655]; 
    assign layer_0[10621] = in[613]; 
    assign layer_0[10622] = in[836] & in[660]; 
    assign layer_0[10623] = ~in[634] | (in[870] & in[634]); 
    assign layer_0[10624] = ~in[791]; 
    assign layer_0[10625] = ~(in[197] & in[855]); 
    assign layer_0[10626] = 1'b1; 
    assign layer_0[10627] = ~(in[140] & in[467]); 
    assign layer_0[10628] = in[250] ^ in[223]; 
    assign layer_0[10629] = ~in[524] | (in[610] & in[524]); 
    assign layer_0[10630] = ~in[603] | (in[603] & in[473]); 
    assign layer_0[10631] = in[894] ^ in[487]; 
    assign layer_0[10632] = ~in[987] | (in[987] & in[465]); 
    assign layer_0[10633] = ~(in[777] | in[721]); 
    assign layer_0[10634] = in[291]; 
    assign layer_0[10635] = ~in[746]; 
    assign layer_0[10636] = ~(in[260] ^ in[452]); 
    assign layer_0[10637] = ~(in[158] ^ in[622]); 
    assign layer_0[10638] = ~in[292]; 
    assign layer_0[10639] = in[932] ^ in[955]; 
    assign layer_0[10640] = in[380] & ~in[886]; 
    assign layer_0[10641] = ~(in[1016] | in[386]); 
    assign layer_0[10642] = ~(in[923] ^ in[681]); 
    assign layer_0[10643] = in[951] ^ in[952]; 
    assign layer_0[10644] = in[368] | in[728]; 
    assign layer_0[10645] = ~(in[676] & in[634]); 
    assign layer_0[10646] = ~in[91] | (in[940] & in[91]); 
    assign layer_0[10647] = ~in[491]; 
    assign layer_0[10648] = ~(in[698] | in[698]); 
    assign layer_0[10649] = ~(in[371] & in[911]); 
    assign layer_0[10650] = in[984] & in[985]; 
    assign layer_0[10651] = ~in[1014]; 
    assign layer_0[10652] = ~(in[937] ^ in[876]); 
    assign layer_0[10653] = ~in[580]; 
    assign layer_0[10654] = ~(in[377] ^ in[451]); 
    assign layer_0[10655] = in[311]; 
    assign layer_0[10656] = ~(in[602] ^ in[523]); 
    assign layer_0[10657] = in[1015] ^ in[747]; 
    assign layer_0[10658] = ~in[68] | (in[68] & in[748]); 
    assign layer_0[10659] = ~(in[583] & in[419]); 
    assign layer_0[10660] = ~(in[522] ^ in[210]); 
    assign layer_0[10661] = in[724] ^ in[460]; 
    assign layer_0[10662] = ~(in[869] ^ in[218]); 
    assign layer_0[10663] = ~(in[578] ^ in[224]); 
    assign layer_0[10664] = in[314] & ~in[938]; 
    assign layer_0[10665] = ~in[451] | (in[451] & in[734]); 
    assign layer_0[10666] = ~in[604] | (in[604] & in[804]); 
    assign layer_0[10667] = in[533] | in[512]; 
    assign layer_0[10668] = ~(in[29] ^ in[259]); 
    assign layer_0[10669] = in[844] ^ in[613]; 
    assign layer_0[10670] = 1'b0; 
    assign layer_0[10671] = ~in[297]; 
    assign layer_0[10672] = ~in[354] | (in[871] & in[354]); 
    assign layer_0[10673] = in[985] & ~in[644]; 
    assign layer_0[10674] = in[327] ^ in[275]; 
    assign layer_0[10675] = ~(in[867] | in[63]); 
    assign layer_0[10676] = ~(in[227] & in[332]); 
    assign layer_0[10677] = ~in[400] | (in[246] & in[400]); 
    assign layer_0[10678] = in[283] ^ in[792]; 
    assign layer_0[10679] = 1'b0; 
    assign layer_0[10680] = in[258] ^ in[463]; 
    assign layer_0[10681] = ~(in[615] ^ in[366]); 
    assign layer_0[10682] = in[978] | in[944]; 
    assign layer_0[10683] = ~(in[692] ^ in[114]); 
    assign layer_0[10684] = in[969]; 
    assign layer_0[10685] = in[129]; 
    assign layer_0[10686] = in[613] & ~in[447]; 
    assign layer_0[10687] = ~(in[809] ^ in[975]); 
    assign layer_0[10688] = in[993] | in[743]; 
    assign layer_0[10689] = ~(in[625] ^ in[195]); 
    assign layer_0[10690] = ~in[147]; 
    assign layer_0[10691] = in[9] ^ in[808]; 
    assign layer_0[10692] = ~(in[708] | in[306]); 
    assign layer_0[10693] = ~in[154]; 
    assign layer_0[10694] = in[183] & ~in[613]; 
    assign layer_0[10695] = in[244] ^ in[97]; 
    assign layer_0[10696] = 1'b0; 
    assign layer_0[10697] = ~(in[504] ^ in[708]); 
    assign layer_0[10698] = in[964] ^ in[265]; 
    assign layer_0[10699] = in[857] ^ in[888]; 
    assign layer_0[10700] = in[999]; 
    assign layer_0[10701] = in[519] ^ in[903]; 
    assign layer_0[10702] = ~(in[11] ^ in[36]); 
    assign layer_0[10703] = 1'b0; 
    assign layer_0[10704] = in[580] | in[763]; 
    assign layer_0[10705] = 1'b1; 
    assign layer_0[10706] = in[550] ^ in[941]; 
    assign layer_0[10707] = ~(in[133] ^ in[295]); 
    assign layer_0[10708] = ~(in[226] & in[932]); 
    assign layer_0[10709] = in[694] ^ in[854]; 
    assign layer_0[10710] = in[603] ^ in[794]; 
    assign layer_0[10711] = in[950] ^ in[725]; 
    assign layer_0[10712] = in[742] & ~in[669]; 
    assign layer_0[10713] = in[655]; 
    assign layer_0[10714] = in[597] ^ in[866]; 
    assign layer_0[10715] = in[248] & in[246]; 
    assign layer_0[10716] = in[799] | in[904]; 
    assign layer_0[10717] = ~(in[727] ^ in[282]); 
    assign layer_0[10718] = in[226] ^ in[596]; 
    assign layer_0[10719] = ~(in[328] | in[684]); 
    assign layer_0[10720] = in[499] & in[423]; 
    assign layer_0[10721] = in[106] & ~in[322]; 
    assign layer_0[10722] = in[958] & ~in[576]; 
    assign layer_0[10723] = ~(in[536] ^ in[872]); 
    assign layer_0[10724] = in[176] ^ in[44]; 
    assign layer_0[10725] = in[276] & ~in[847]; 
    assign layer_0[10726] = in[24] | in[959]; 
    assign layer_0[10727] = ~(in[918] ^ in[519]); 
    assign layer_0[10728] = in[857] | in[383]; 
    assign layer_0[10729] = in[527]; 
    assign layer_0[10730] = in[372] & ~in[904]; 
    assign layer_0[10731] = in[332] ^ in[716]; 
    assign layer_0[10732] = ~(in[245] ^ in[316]); 
    assign layer_0[10733] = ~in[874]; 
    assign layer_0[10734] = 1'b0; 
    assign layer_0[10735] = in[766] ^ in[344]; 
    assign layer_0[10736] = ~(in[237] & in[755]); 
    assign layer_0[10737] = in[508] ^ in[174]; 
    assign layer_0[10738] = ~(in[724] | in[3]); 
    assign layer_0[10739] = ~in[821] | (in[285] & in[821]); 
    assign layer_0[10740] = ~in[473] | (in[473] & in[66]); 
    assign layer_0[10741] = ~(in[596] | in[489]); 
    assign layer_0[10742] = in[85] & ~in[933]; 
    assign layer_0[10743] = in[294] ^ in[194]; 
    assign layer_0[10744] = in[251] & in[56]; 
    assign layer_0[10745] = ~(in[916] | in[900]); 
    assign layer_0[10746] = ~(in[3] ^ in[51]); 
    assign layer_0[10747] = ~(in[905] ^ in[904]); 
    assign layer_0[10748] = ~in[66] | (in[66] & in[837]); 
    assign layer_0[10749] = in[920] & in[162]; 
    assign layer_0[10750] = ~(in[505] ^ in[379]); 
    assign layer_0[10751] = in[955] & ~in[929]; 
    assign layer_0[10752] = in[659] & ~in[955]; 
    assign layer_0[10753] = 1'b0; 
    assign layer_0[10754] = ~in[568] | (in[858] & in[568]); 
    assign layer_0[10755] = in[563] & in[157]; 
    assign layer_0[10756] = ~(in[619] ^ in[789]); 
    assign layer_0[10757] = in[910] ^ in[583]; 
    assign layer_0[10758] = ~in[628]; 
    assign layer_0[10759] = in[466]; 
    assign layer_0[10760] = in[628] & ~in[827]; 
    assign layer_0[10761] = ~(in[985] & in[540]); 
    assign layer_0[10762] = ~(in[89] ^ in[825]); 
    assign layer_0[10763] = ~(in[873] ^ in[904]); 
    assign layer_0[10764] = in[761] | in[860]; 
    assign layer_0[10765] = ~(in[982] ^ in[745]); 
    assign layer_0[10766] = ~(in[809] ^ in[836]); 
    assign layer_0[10767] = in[458] ^ in[840]; 
    assign layer_0[10768] = ~(in[260] ^ in[450]); 
    assign layer_0[10769] = ~in[121]; 
    assign layer_0[10770] = in[475] & in[473]; 
    assign layer_0[10771] = in[871] & ~in[652]; 
    assign layer_0[10772] = ~in[756] | (in[756] & in[414]); 
    assign layer_0[10773] = 1'b1; 
    assign layer_0[10774] = ~(in[322] ^ in[508]); 
    assign layer_0[10775] = in[489] & ~in[243]; 
    assign layer_0[10776] = ~in[843]; 
    assign layer_0[10777] = ~(in[683] & in[46]); 
    assign layer_0[10778] = in[520] ^ in[200]; 
    assign layer_0[10779] = in[934] & ~in[384]; 
    assign layer_0[10780] = ~(in[779] | in[523]); 
    assign layer_0[10781] = in[671]; 
    assign layer_0[10782] = ~in[568]; 
    assign layer_0[10783] = in[744]; 
    assign layer_0[10784] = ~(in[338] ^ in[175]); 
    assign layer_0[10785] = ~in[91]; 
    assign layer_0[10786] = in[279] & ~in[550]; 
    assign layer_0[10787] = in[143] ^ in[365]; 
    assign layer_0[10788] = ~(in[984] ^ in[490]); 
    assign layer_0[10789] = in[756] | in[627]; 
    assign layer_0[10790] = ~in[493]; 
    assign layer_0[10791] = ~in[735]; 
    assign layer_0[10792] = ~(in[222] ^ in[555]); 
    assign layer_0[10793] = in[919] & ~in[810]; 
    assign layer_0[10794] = in[604]; 
    assign layer_0[10795] = in[396] ^ in[492]; 
    assign layer_0[10796] = ~in[522]; 
    assign layer_0[10797] = in[657] ^ in[970]; 
    assign layer_0[10798] = in[346] ^ in[968]; 
    assign layer_0[10799] = in[751] | in[835]; 
    assign layer_0[10800] = ~in[358] | (in[358] & in[300]); 
    assign layer_0[10801] = ~in[145] | (in[145] & in[176]); 
    assign layer_0[10802] = ~(in[467] ^ in[681]); 
    assign layer_0[10803] = ~(in[603] & in[342]); 
    assign layer_0[10804] = ~(in[974] | in[111]); 
    assign layer_0[10805] = in[319] ^ in[688]; 
    assign layer_0[10806] = ~in[260]; 
    assign layer_0[10807] = ~(in[437] ^ in[221]); 
    assign layer_0[10808] = in[343] ^ in[309]; 
    assign layer_0[10809] = in[465] & ~in[773]; 
    assign layer_0[10810] = in[79] & ~in[42]; 
    assign layer_0[10811] = ~in[823] | (in[847] & in[823]); 
    assign layer_0[10812] = in[77] & ~in[260]; 
    assign layer_0[10813] = ~(in[500] ^ in[759]); 
    assign layer_0[10814] = in[153] & ~in[740]; 
    assign layer_0[10815] = ~in[772]; 
    assign layer_0[10816] = ~(in[915] ^ in[543]); 
    assign layer_0[10817] = in[887]; 
    assign layer_0[10818] = ~(in[822] ^ in[917]); 
    assign layer_0[10819] = ~(in[840] ^ in[498]); 
    assign layer_0[10820] = in[269] & ~in[1016]; 
    assign layer_0[10821] = in[900]; 
    assign layer_0[10822] = in[481] & in[535]; 
    assign layer_0[10823] = in[569] ^ in[536]; 
    assign layer_0[10824] = in[238] ^ in[262]; 
    assign layer_0[10825] = in[609] | in[379]; 
    assign layer_0[10826] = in[458] & ~in[268]; 
    assign layer_0[10827] = in[466] ^ in[655]; 
    assign layer_0[10828] = ~in[533] | (in[533] & in[861]); 
    assign layer_0[10829] = ~(in[504] ^ in[871]); 
    assign layer_0[10830] = in[134]; 
    assign layer_0[10831] = ~in[937]; 
    assign layer_0[10832] = in[1014]; 
    assign layer_0[10833] = ~in[884]; 
    assign layer_0[10834] = in[594]; 
    assign layer_0[10835] = in[347] & in[1015]; 
    assign layer_0[10836] = ~(in[533] ^ in[414]); 
    assign layer_0[10837] = ~in[117] | (in[117] & in[771]); 
    assign layer_0[10838] = ~in[357] | (in[357] & in[878]); 
    assign layer_0[10839] = ~(in[730] ^ in[538]); 
    assign layer_0[10840] = in[573] ^ in[788]; 
    assign layer_0[10841] = in[28] ^ in[533]; 
    assign layer_0[10842] = ~in[889] | (in[790] & in[889]); 
    assign layer_0[10843] = ~(in[264] ^ in[732]); 
    assign layer_0[10844] = in[110] ^ in[922]; 
    assign layer_0[10845] = ~in[872]; 
    assign layer_0[10846] = ~(in[341] ^ in[935]); 
    assign layer_0[10847] = ~in[81] | (in[533] & in[81]); 
    assign layer_0[10848] = in[536]; 
    assign layer_0[10849] = in[420] & ~in[46]; 
    assign layer_0[10850] = ~in[869]; 
    assign layer_0[10851] = in[249] | in[510]; 
    assign layer_0[10852] = in[522] | in[97]; 
    assign layer_0[10853] = in[477] | in[918]; 
    assign layer_0[10854] = ~(in[1021] ^ in[491]); 
    assign layer_0[10855] = ~in[582] | (in[904] & in[582]); 
    assign layer_0[10856] = in[85] ^ in[1017]; 
    assign layer_0[10857] = in[707]; 
    assign layer_0[10858] = ~in[60]; 
    assign layer_0[10859] = ~(in[840] ^ in[887]); 
    assign layer_0[10860] = ~in[650] | (in[650] & in[238]); 
    assign layer_0[10861] = in[179]; 
    assign layer_0[10862] = in[853] ^ in[657]; 
    assign layer_0[10863] = in[110] ^ in[261]; 
    assign layer_0[10864] = ~in[867]; 
    assign layer_0[10865] = in[982]; 
    assign layer_0[10866] = ~(in[931] ^ in[325]); 
    assign layer_0[10867] = ~in[311]; 
    assign layer_0[10868] = ~(in[810] ^ in[246]); 
    assign layer_0[10869] = ~in[407]; 
    assign layer_0[10870] = ~(in[12] ^ in[485]); 
    assign layer_0[10871] = in[601] ^ in[935]; 
    assign layer_0[10872] = in[12] & ~in[81]; 
    assign layer_0[10873] = ~in[77] | (in[657] & in[77]); 
    assign layer_0[10874] = ~in[737]; 
    assign layer_0[10875] = ~(in[618] & in[474]); 
    assign layer_0[10876] = ~(in[1001] | in[362]); 
    assign layer_0[10877] = in[145] & ~in[796]; 
    assign layer_0[10878] = in[837]; 
    assign layer_0[10879] = ~(in[261] ^ in[177]); 
    assign layer_0[10880] = in[279] ^ in[293]; 
    assign layer_0[10881] = ~in[624]; 
    assign layer_0[10882] = in[994] ^ in[856]; 
    assign layer_0[10883] = in[383]; 
    assign layer_0[10884] = ~(in[472] & in[184]); 
    assign layer_0[10885] = ~(in[888] ^ in[857]); 
    assign layer_0[10886] = 1'b0; 
    assign layer_0[10887] = in[910] | in[567]; 
    assign layer_0[10888] = in[49] & in[302]; 
    assign layer_0[10889] = ~(in[193] & in[689]); 
    assign layer_0[10890] = 1'b0; 
    assign layer_0[10891] = ~in[588] | (in[551] & in[588]); 
    assign layer_0[10892] = ~(in[773] | in[661]); 
    assign layer_0[10893] = ~in[369] | (in[369] & in[885]); 
    assign layer_0[10894] = in[568] ^ in[300]; 
    assign layer_0[10895] = ~(in[936] ^ in[968]); 
    assign layer_0[10896] = in[621] ^ in[492]; 
    assign layer_0[10897] = in[643] | in[520]; 
    assign layer_0[10898] = in[59] ^ in[774]; 
    assign layer_0[10899] = in[182] & ~in[713]; 
    assign layer_0[10900] = 1'b0; 
    assign layer_0[10901] = in[611] ^ in[110]; 
    assign layer_0[10902] = ~in[119] | (in[534] & in[119]); 
    assign layer_0[10903] = ~(in[239] | in[778]); 
    assign layer_0[10904] = ~in[844] | (in[844] & in[947]); 
    assign layer_0[10905] = ~(in[276] ^ in[461]); 
    assign layer_0[10906] = in[80] ^ in[937]; 
    assign layer_0[10907] = ~in[666] | (in[996] & in[666]); 
    assign layer_0[10908] = in[521] ^ in[824]; 
    assign layer_0[10909] = ~(in[707] ^ in[97]); 
    assign layer_0[10910] = ~(in[299] ^ in[839]); 
    assign layer_0[10911] = ~(in[264] ^ in[660]); 
    assign layer_0[10912] = ~(in[174] ^ in[643]); 
    assign layer_0[10913] = ~(in[717] & in[601]); 
    assign layer_0[10914] = in[437] & ~in[848]; 
    assign layer_0[10915] = in[352] | in[386]; 
    assign layer_0[10916] = ~(in[328] & in[478]); 
    assign layer_0[10917] = in[641]; 
    assign layer_0[10918] = ~(in[210] ^ in[635]); 
    assign layer_0[10919] = ~(in[284] | in[403]); 
    assign layer_0[10920] = in[614] & ~in[531]; 
    assign layer_0[10921] = in[736]; 
    assign layer_0[10922] = in[50] ^ in[531]; 
    assign layer_0[10923] = in[50] ^ in[467]; 
    assign layer_0[10924] = ~(in[757] ^ in[747]); 
    assign layer_0[10925] = in[904]; 
    assign layer_0[10926] = in[67]; 
    assign layer_0[10927] = 1'b1; 
    assign layer_0[10928] = in[821] ^ in[854]; 
    assign layer_0[10929] = ~in[601] | (in[601] & in[809]); 
    assign layer_0[10930] = ~in[714] | (in[249] & in[714]); 
    assign layer_0[10931] = ~in[504] | (in[939] & in[504]); 
    assign layer_0[10932] = ~in[984] | (in[890] & in[984]); 
    assign layer_0[10933] = ~in[795]; 
    assign layer_0[10934] = in[905]; 
    assign layer_0[10935] = in[508] & in[998]; 
    assign layer_0[10936] = in[206] ^ in[588]; 
    assign layer_0[10937] = ~(in[267] | in[622]); 
    assign layer_0[10938] = in[489] ^ in[224]; 
    assign layer_0[10939] = ~in[862] | (in[779] & in[862]); 
    assign layer_0[10940] = ~in[836] | (in[836] & in[509]); 
    assign layer_0[10941] = in[475] ^ in[442]; 
    assign layer_0[10942] = ~(in[77] | in[33]); 
    assign layer_0[10943] = ~in[452]; 
    assign layer_0[10944] = in[646] & ~in[538]; 
    assign layer_0[10945] = 1'b0; 
    assign layer_0[10946] = in[709] & ~in[679]; 
    assign layer_0[10947] = ~(in[28] & in[500]); 
    assign layer_0[10948] = ~in[838] | (in[717] & in[838]); 
    assign layer_0[10949] = in[964] ^ in[588]; 
    assign layer_0[10950] = in[468] ^ in[616]; 
    assign layer_0[10951] = ~(in[360] & in[695]); 
    assign layer_0[10952] = ~(in[98] ^ in[665]); 
    assign layer_0[10953] = ~(in[644] | in[556]); 
    assign layer_0[10954] = in[451] & ~in[626]; 
    assign layer_0[10955] = ~(in[905] ^ in[760]); 
    assign layer_0[10956] = in[126] | in[409]; 
    assign layer_0[10957] = in[161] ^ in[314]; 
    assign layer_0[10958] = in[603] ^ in[843]; 
    assign layer_0[10959] = in[760]; 
    assign layer_0[10960] = in[301]; 
    assign layer_0[10961] = ~(in[901] ^ in[688]); 
    assign layer_0[10962] = ~(in[574] | in[680]); 
    assign layer_0[10963] = ~(in[715] ^ in[701]); 
    assign layer_0[10964] = ~in[789]; 
    assign layer_0[10965] = in[868] & in[908]; 
    assign layer_0[10966] = in[284]; 
    assign layer_0[10967] = in[831] | in[907]; 
    assign layer_0[10968] = in[607] & ~in[116]; 
    assign layer_0[10969] = ~in[195]; 
    assign layer_0[10970] = ~in[987]; 
    assign layer_0[10971] = in[966]; 
    assign layer_0[10972] = ~(in[111] ^ in[1006]); 
    assign layer_0[10973] = in[604] ^ in[278]; 
    assign layer_0[10974] = ~in[261] | (in[580] & in[261]); 
    assign layer_0[10975] = in[206]; 
    assign layer_0[10976] = 1'b1; 
    assign layer_0[10977] = in[717] & ~in[945]; 
    assign layer_0[10978] = 1'b0; 
    assign layer_0[10979] = in[878]; 
    assign layer_0[10980] = in[317] ^ in[904]; 
    assign layer_0[10981] = in[981] & ~in[916]; 
    assign layer_0[10982] = ~(in[948] | in[940]); 
    assign layer_0[10983] = in[519] & ~in[465]; 
    assign layer_0[10984] = ~in[701] | (in[38] & in[701]); 
    assign layer_0[10985] = ~in[575]; 
    assign layer_0[10986] = in[424] & in[161]; 
    assign layer_0[10987] = in[444] ^ in[825]; 
    assign layer_0[10988] = in[854] ^ in[691]; 
    assign layer_0[10989] = in[623] ^ in[714]; 
    assign layer_0[10990] = in[294] | in[645]; 
    assign layer_0[10991] = in[761] & ~in[915]; 
    assign layer_0[10992] = ~(in[286] | in[701]); 
    assign layer_0[10993] = ~(in[684] ^ in[916]); 
    assign layer_0[10994] = ~in[716] | (in[716] & in[7]); 
    assign layer_0[10995] = ~in[58] | (in[313] & in[58]); 
    assign layer_0[10996] = in[535] & in[635]; 
    assign layer_0[10997] = ~(in[866] | in[757]); 
    assign layer_0[10998] = in[618]; 
    assign layer_0[10999] = ~(in[511] & in[781]); 
    assign layer_0[11000] = in[239]; 
    assign layer_0[11001] = ~(in[889] ^ in[969]); 
    assign layer_0[11002] = ~in[437] | (in[590] & in[437]); 
    assign layer_0[11003] = in[584]; 
    assign layer_0[11004] = ~in[885] | (in[885] & in[883]); 
    assign layer_0[11005] = ~in[347] | (in[748] & in[347]); 
    assign layer_0[11006] = ~(in[300] | in[348]); 
    assign layer_0[11007] = ~(in[679] & in[599]); 
    assign layer_0[11008] = 1'b1; 
    assign layer_0[11009] = ~(in[775] | in[980]); 
    assign layer_0[11010] = ~in[536]; 
    assign layer_0[11011] = ~(in[523] ^ in[280]); 
    assign layer_0[11012] = in[843] ^ in[859]; 
    assign layer_0[11013] = in[187] | in[91]; 
    assign layer_0[11014] = ~(in[948] | in[1003]); 
    assign layer_0[11015] = ~(in[60] ^ in[12]); 
    assign layer_0[11016] = in[807] ^ in[264]; 
    assign layer_0[11017] = ~(in[13] | in[1013]); 
    assign layer_0[11018] = ~in[875]; 
    assign layer_0[11019] = in[113] ^ in[7]; 
    assign layer_0[11020] = ~(in[521] ^ in[572]); 
    assign layer_0[11021] = ~in[379]; 
    assign layer_0[11022] = in[648] & ~in[350]; 
    assign layer_0[11023] = ~in[598]; 
    assign layer_0[11024] = ~(in[522] ^ in[510]); 
    assign layer_0[11025] = ~in[829]; 
    assign layer_0[11026] = in[914] ^ in[978]; 
    assign layer_0[11027] = in[791] ^ in[505]; 
    assign layer_0[11028] = in[585] ^ in[566]; 
    assign layer_0[11029] = ~in[348]; 
    assign layer_0[11030] = ~in[153] | (in[153] & in[499]); 
    assign layer_0[11031] = ~(in[125] | in[938]); 
    assign layer_0[11032] = in[127] & ~in[533]; 
    assign layer_0[11033] = ~(in[748] | in[353]); 
    assign layer_0[11034] = ~(in[607] ^ in[658]); 
    assign layer_0[11035] = ~(in[515] | in[886]); 
    assign layer_0[11036] = in[687]; 
    assign layer_0[11037] = in[627]; 
    assign layer_0[11038] = in[828] ^ in[494]; 
    assign layer_0[11039] = ~(in[820] | in[556]); 
    assign layer_0[11040] = in[916]; 
    assign layer_0[11041] = in[31] & ~in[809]; 
    assign layer_0[11042] = ~(in[827] ^ in[350]); 
    assign layer_0[11043] = ~in[52] | (in[52] & in[557]); 
    assign layer_0[11044] = ~in[670] | (in[829] & in[670]); 
    assign layer_0[11045] = ~in[140] | (in[140] & in[748]); 
    assign layer_0[11046] = ~in[852] | (in[852] & in[907]); 
    assign layer_0[11047] = ~(in[337] ^ in[483]); 
    assign layer_0[11048] = ~in[870] | (in[870] & in[477]); 
    assign layer_0[11049] = ~(in[955] ^ in[886]); 
    assign layer_0[11050] = ~in[412] | (in[521] & in[412]); 
    assign layer_0[11051] = ~(in[23] ^ in[894]); 
    assign layer_0[11052] = in[883] | in[990]; 
    assign layer_0[11053] = ~in[141]; 
    assign layer_0[11054] = ~in[412]; 
    assign layer_0[11055] = ~in[870] | (in[870] & in[918]); 
    assign layer_0[11056] = in[0]; 
    assign layer_0[11057] = in[875] ^ in[955]; 
    assign layer_0[11058] = in[646] ^ in[220]; 
    assign layer_0[11059] = in[189]; 
    assign layer_0[11060] = in[119] & in[534]; 
    assign layer_0[11061] = ~in[300] | (in[834] & in[300]); 
    assign layer_0[11062] = ~in[397] | (in[683] & in[397]); 
    assign layer_0[11063] = ~(in[599] | in[317]); 
    assign layer_0[11064] = ~in[281] | (in[17] & in[281]); 
    assign layer_0[11065] = in[984] & ~in[603]; 
    assign layer_0[11066] = in[259] & ~in[331]; 
    assign layer_0[11067] = in[762] ^ in[984]; 
    assign layer_0[11068] = ~(in[145] & in[421]); 
    assign layer_0[11069] = in[572] | in[266]; 
    assign layer_0[11070] = ~in[205]; 
    assign layer_0[11071] = ~(in[699] ^ in[659]); 
    assign layer_0[11072] = ~in[96]; 
    assign layer_0[11073] = ~(in[900] ^ in[841]); 
    assign layer_0[11074] = ~in[6]; 
    assign layer_0[11075] = in[449] & ~in[260]; 
    assign layer_0[11076] = in[449] | in[949]; 
    assign layer_0[11077] = ~(in[922] ^ in[220]); 
    assign layer_0[11078] = ~(in[622] | in[808]); 
    assign layer_0[11079] = in[218] ^ in[746]; 
    assign layer_0[11080] = in[309] ^ in[851]; 
    assign layer_0[11081] = ~(in[544] & in[739]); 
    assign layer_0[11082] = in[117] ^ in[155]; 
    assign layer_0[11083] = ~(in[949] ^ in[307]); 
    assign layer_0[11084] = ~in[911]; 
    assign layer_0[11085] = ~(in[319] & in[840]); 
    assign layer_0[11086] = in[130] & in[337]; 
    assign layer_0[11087] = in[810] | in[651]; 
    assign layer_0[11088] = ~in[811]; 
    assign layer_0[11089] = in[535] | in[800]; 
    assign layer_0[11090] = ~(in[762] ^ in[757]); 
    assign layer_0[11091] = in[810] & in[45]; 
    assign layer_0[11092] = in[289] & ~in[203]; 
    assign layer_0[11093] = ~(in[981] ^ in[982]); 
    assign layer_0[11094] = ~in[97]; 
    assign layer_0[11095] = ~(in[68] & in[419]); 
    assign layer_0[11096] = ~(in[732] ^ in[749]); 
    assign layer_0[11097] = in[361] ^ in[965]; 
    assign layer_0[11098] = in[436] ^ in[716]; 
    assign layer_0[11099] = in[182] & in[460]; 
    assign layer_0[11100] = in[224] | in[762]; 
    assign layer_0[11101] = in[584] & ~in[830]; 
    assign layer_0[11102] = ~in[434]; 
    assign layer_0[11103] = ~in[584] | (in[986] & in[584]); 
    assign layer_0[11104] = ~in[539]; 
    assign layer_0[11105] = in[396] & ~in[224]; 
    assign layer_0[11106] = in[354] | in[291]; 
    assign layer_0[11107] = ~(in[653] | in[136]); 
    assign layer_0[11108] = in[785] & ~in[401]; 
    assign layer_0[11109] = ~(in[399] ^ in[970]); 
    assign layer_0[11110] = in[397] & ~in[588]; 
    assign layer_0[11111] = in[832] | in[359]; 
    assign layer_0[11112] = in[117]; 
    assign layer_0[11113] = in[856] & ~in[855]; 
    assign layer_0[11114] = ~in[264]; 
    assign layer_0[11115] = ~(in[266] ^ in[835]); 
    assign layer_0[11116] = in[358] | in[633]; 
    assign layer_0[11117] = in[857] | in[349]; 
    assign layer_0[11118] = in[1020]; 
    assign layer_0[11119] = in[665] ^ in[676]; 
    assign layer_0[11120] = ~in[648] | (in[868] & in[648]); 
    assign layer_0[11121] = in[986] ^ in[757]; 
    assign layer_0[11122] = ~(in[955] ^ in[889]); 
    assign layer_0[11123] = in[940]; 
    assign layer_0[11124] = in[622] & ~in[919]; 
    assign layer_0[11125] = in[491]; 
    assign layer_0[11126] = in[552] ^ in[483]; 
    assign layer_0[11127] = ~(in[261] ^ in[285]); 
    assign layer_0[11128] = in[535] & ~in[662]; 
    assign layer_0[11129] = in[857]; 
    assign layer_0[11130] = in[256] | in[96]; 
    assign layer_0[11131] = ~in[238]; 
    assign layer_0[11132] = in[963] & ~in[950]; 
    assign layer_0[11133] = in[572] ^ in[505]; 
    assign layer_0[11134] = ~(in[1017] ^ in[149]); 
    assign layer_0[11135] = in[250] | in[865]; 
    assign layer_0[11136] = ~in[860] | (in[860] & in[855]); 
    assign layer_0[11137] = ~in[906]; 
    assign layer_0[11138] = ~(in[887] ^ in[884]); 
    assign layer_0[11139] = ~in[588] | (in[286] & in[588]); 
    assign layer_0[11140] = in[918] ^ in[970]; 
    assign layer_0[11141] = in[812]; 
    assign layer_0[11142] = in[923] ^ in[343]; 
    assign layer_0[11143] = ~(in[335] ^ in[716]); 
    assign layer_0[11144] = in[34]; 
    assign layer_0[11145] = ~(in[983] ^ in[967]); 
    assign layer_0[11146] = ~(in[635] | in[756]); 
    assign layer_0[11147] = in[858] ^ in[856]; 
    assign layer_0[11148] = ~(in[791] & in[937]); 
    assign layer_0[11149] = in[657] ^ in[73]; 
    assign layer_0[11150] = ~(in[501] ^ in[405]); 
    assign layer_0[11151] = in[411] | in[48]; 
    assign layer_0[11152] = ~in[744]; 
    assign layer_0[11153] = in[194] ^ in[261]; 
    assign layer_0[11154] = ~in[73] | (in[73] & in[108]); 
    assign layer_0[11155] = in[967] & ~in[837]; 
    assign layer_0[11156] = ~(in[958] & in[784]); 
    assign layer_0[11157] = in[591] & ~in[572]; 
    assign layer_0[11158] = ~(in[492] | in[127]); 
    assign layer_0[11159] = ~in[148]; 
    assign layer_0[11160] = ~(in[919] & in[631]); 
    assign layer_0[11161] = ~in[55]; 
    assign layer_0[11162] = ~in[1016]; 
    assign layer_0[11163] = in[789] ^ in[618]; 
    assign layer_0[11164] = ~in[734] | (in[734] & in[745]); 
    assign layer_0[11165] = in[468] | in[982]; 
    assign layer_0[11166] = ~(in[56] ^ in[656]); 
    assign layer_0[11167] = in[759] ^ in[565]; 
    assign layer_0[11168] = in[787] ^ in[477]; 
    assign layer_0[11169] = ~in[667] | (in[667] & in[177]); 
    assign layer_0[11170] = ~(in[622] ^ in[655]); 
    assign layer_0[11171] = in[179] & ~in[435]; 
    assign layer_0[11172] = ~in[329]; 
    assign layer_0[11173] = in[699] | in[902]; 
    assign layer_0[11174] = ~(in[438] & in[249]); 
    assign layer_0[11175] = ~(in[935] ^ in[966]); 
    assign layer_0[11176] = in[839]; 
    assign layer_0[11177] = in[1004] ^ in[331]; 
    assign layer_0[11178] = ~in[350] | (in[351] & in[350]); 
    assign layer_0[11179] = in[854] ^ in[354]; 
    assign layer_0[11180] = ~in[900]; 
    assign layer_0[11181] = in[339] | in[348]; 
    assign layer_0[11182] = in[809] ^ in[573]; 
    assign layer_0[11183] = in[337]; 
    assign layer_0[11184] = ~(in[989] ^ in[932]); 
    assign layer_0[11185] = ~(in[48] ^ in[508]); 
    assign layer_0[11186] = in[262] & ~in[823]; 
    assign layer_0[11187] = in[370] | in[223]; 
    assign layer_0[11188] = in[189] | in[912]; 
    assign layer_0[11189] = ~(in[537] | in[741]); 
    assign layer_0[11190] = in[940] ^ in[275]; 
    assign layer_0[11191] = in[541]; 
    assign layer_0[11192] = ~in[1020]; 
    assign layer_0[11193] = in[311] & in[396]; 
    assign layer_0[11194] = ~in[17]; 
    assign layer_0[11195] = ~(in[1000] | in[605]); 
    assign layer_0[11196] = ~in[291]; 
    assign layer_0[11197] = in[19] & in[483]; 
    assign layer_0[11198] = ~(in[823] ^ in[855]); 
    assign layer_0[11199] = ~in[714] | (in[714] & in[949]); 
    assign layer_0[11200] = in[92] & in[260]; 
    assign layer_0[11201] = ~(in[102] ^ in[584]); 
    assign layer_0[11202] = in[660] & in[365]; 
    assign layer_0[11203] = in[828] ^ in[693]; 
    assign layer_0[11204] = ~in[707]; 
    assign layer_0[11205] = in[650] & ~in[30]; 
    assign layer_0[11206] = ~in[899]; 
    assign layer_0[11207] = in[518] ^ in[50]; 
    assign layer_0[11208] = in[3]; 
    assign layer_0[11209] = in[75] & ~in[145]; 
    assign layer_0[11210] = in[836] | in[463]; 
    assign layer_0[11211] = ~(in[18] ^ in[876]); 
    assign layer_0[11212] = in[707] ^ in[302]; 
    assign layer_0[11213] = ~(in[11] ^ in[661]); 
    assign layer_0[11214] = in[888] & ~in[889]; 
    assign layer_0[11215] = in[203]; 
    assign layer_0[11216] = in[267] ^ in[648]; 
    assign layer_0[11217] = ~in[373] | (in[373] & in[1015]); 
    assign layer_0[11218] = in[426]; 
    assign layer_0[11219] = ~(in[94] ^ in[750]); 
    assign layer_0[11220] = ~in[380] | (in[380] & in[159]); 
    assign layer_0[11221] = in[969] ^ in[968]; 
    assign layer_0[11222] = ~(in[268] ^ in[67]); 
    assign layer_0[11223] = in[484] ^ in[597]; 
    assign layer_0[11224] = ~in[40] | (in[260] & in[40]); 
    assign layer_0[11225] = in[265] ^ in[262]; 
    assign layer_0[11226] = in[492] & ~in[616]; 
    assign layer_0[11227] = in[981] & ~in[827]; 
    assign layer_0[11228] = in[378] & ~in[1016]; 
    assign layer_0[11229] = ~in[194] | (in[299] & in[194]); 
    assign layer_0[11230] = in[112] ^ in[687]; 
    assign layer_0[11231] = ~(in[640] ^ in[343]); 
    assign layer_0[11232] = ~(in[612] ^ in[402]); 
    assign layer_0[11233] = in[937] | in[936]; 
    assign layer_0[11234] = ~(in[364] ^ in[48]); 
    assign layer_0[11235] = in[44] | in[588]; 
    assign layer_0[11236] = ~(in[692] & in[416]); 
    assign layer_0[11237] = ~in[763]; 
    assign layer_0[11238] = ~in[467] | (in[715] & in[467]); 
    assign layer_0[11239] = ~(in[506] ^ in[645]); 
    assign layer_0[11240] = ~(in[547] ^ in[608]); 
    assign layer_0[11241] = in[573]; 
    assign layer_0[11242] = in[324] ^ in[967]; 
    assign layer_0[11243] = ~in[18]; 
    assign layer_0[11244] = ~(in[885] ^ in[883]); 
    assign layer_0[11245] = in[635] & in[329]; 
    assign layer_0[11246] = in[858] | in[937]; 
    assign layer_0[11247] = ~in[997] | (in[997] & in[986]); 
    assign layer_0[11248] = ~(in[148] & in[825]); 
    assign layer_0[11249] = ~(in[650] ^ in[660]); 
    assign layer_0[11250] = ~(in[19] ^ in[937]); 
    assign layer_0[11251] = ~in[634] | (in[917] & in[634]); 
    assign layer_0[11252] = ~in[428] | (in[857] & in[428]); 
    assign layer_0[11253] = in[880] | in[364]; 
    assign layer_0[11254] = in[611] | in[852]; 
    assign layer_0[11255] = in[566] & ~in[652]; 
    assign layer_0[11256] = ~in[991]; 
    assign layer_0[11257] = ~(in[113] | in[115]); 
    assign layer_0[11258] = ~in[549]; 
    assign layer_0[11259] = ~(in[611] ^ in[645]); 
    assign layer_0[11260] = ~in[433] | (in[433] & in[534]); 
    assign layer_0[11261] = in[489]; 
    assign layer_0[11262] = ~in[324] | (in[324] & in[613]); 
    assign layer_0[11263] = in[617] ^ in[969]; 
    assign layer_0[11264] = ~(in[368] ^ in[955]); 
    assign layer_0[11265] = ~in[791] | (in[791] & in[810]); 
    assign layer_0[11266] = in[84]; 
    assign layer_0[11267] = ~(in[602] ^ in[680]); 
    assign layer_0[11268] = in[843] & in[580]; 
    assign layer_0[11269] = ~(in[455] & in[163]); 
    assign layer_0[11270] = ~in[634]; 
    assign layer_0[11271] = in[128] & ~in[972]; 
    assign layer_0[11272] = ~(in[993] ^ in[599]); 
    assign layer_0[11273] = ~in[147] | (in[918] & in[147]); 
    assign layer_0[11274] = ~(in[123] ^ in[486]); 
    assign layer_0[11275] = in[22]; 
    assign layer_0[11276] = in[490] ^ in[843]; 
    assign layer_0[11277] = ~(in[86] & in[869]); 
    assign layer_0[11278] = in[540] | in[354]; 
    assign layer_0[11279] = in[552] & in[362]; 
    assign layer_0[11280] = ~in[84]; 
    assign layer_0[11281] = in[685] ^ in[122]; 
    assign layer_0[11282] = ~(in[595] | in[6]); 
    assign layer_0[11283] = ~in[389]; 
    assign layer_0[11284] = ~(in[867] ^ in[283]); 
    assign layer_0[11285] = ~(in[925] | in[364]); 
    assign layer_0[11286] = in[376]; 
    assign layer_0[11287] = ~(in[226] ^ in[292]); 
    assign layer_0[11288] = ~in[566]; 
    assign layer_0[11289] = ~(in[481] | in[335]); 
    assign layer_0[11290] = in[446] & in[462]; 
    assign layer_0[11291] = in[233] & ~in[252]; 
    assign layer_0[11292] = ~(in[765] ^ in[873]); 
    assign layer_0[11293] = ~(in[665] ^ in[1004]); 
    assign layer_0[11294] = ~in[874]; 
    assign layer_0[11295] = ~(in[970] ^ in[827]); 
    assign layer_0[11296] = in[133] & in[682]; 
    assign layer_0[11297] = ~in[952]; 
    assign layer_0[11298] = ~(in[628] ^ in[689]); 
    assign layer_0[11299] = in[713] & ~in[637]; 
    assign layer_0[11300] = in[352] ^ in[34]; 
    assign layer_0[11301] = in[434] & in[320]; 
    assign layer_0[11302] = in[899] & in[427]; 
    assign layer_0[11303] = in[555] & ~in[844]; 
    assign layer_0[11304] = ~in[108]; 
    assign layer_0[11305] = ~(in[901] ^ in[950]); 
    assign layer_0[11306] = in[338]; 
    assign layer_0[11307] = ~in[865]; 
    assign layer_0[11308] = ~(in[838] ^ in[937]); 
    assign layer_0[11309] = 1'b0; 
    assign layer_0[11310] = ~(in[984] ^ in[835]); 
    assign layer_0[11311] = in[584]; 
    assign layer_0[11312] = ~(in[569] ^ in[284]); 
    assign layer_0[11313] = ~(in[7] | in[865]); 
    assign layer_0[11314] = in[221] ^ in[854]; 
    assign layer_0[11315] = ~(in[735] ^ in[894]); 
    assign layer_0[11316] = in[910] & in[894]; 
    assign layer_0[11317] = ~(in[324] ^ in[877]); 
    assign layer_0[11318] = in[1002] | in[577]; 
    assign layer_0[11319] = in[824] & ~in[920]; 
    assign layer_0[11320] = ~in[667]; 
    assign layer_0[11321] = in[285] ^ in[903]; 
    assign layer_0[11322] = ~in[370] | (in[707] & in[370]); 
    assign layer_0[11323] = ~(in[732] ^ in[245]); 
    assign layer_0[11324] = in[640]; 
    assign layer_0[11325] = 1'b1; 
    assign layer_0[11326] = ~(in[704] ^ in[219]); 
    assign layer_0[11327] = in[476] & ~in[253]; 
    assign layer_0[11328] = in[195]; 
    assign layer_0[11329] = ~in[146] | (in[622] & in[146]); 
    assign layer_0[11330] = ~(in[827] ^ in[651]); 
    assign layer_0[11331] = in[1013] | in[629]; 
    assign layer_0[11332] = ~in[288]; 
    assign layer_0[11333] = in[676] | in[789]; 
    assign layer_0[11334] = in[952] & in[585]; 
    assign layer_0[11335] = ~(in[954] | in[908]); 
    assign layer_0[11336] = ~(in[519] & in[743]); 
    assign layer_0[11337] = ~(in[254] ^ in[652]); 
    assign layer_0[11338] = ~(in[872] ^ in[844]); 
    assign layer_0[11339] = ~in[648] | (in[557] & in[648]); 
    assign layer_0[11340] = in[508] ^ in[267]; 
    assign layer_0[11341] = in[672]; 
    assign layer_0[11342] = 1'b0; 
    assign layer_0[11343] = ~in[645] | (in[871] & in[645]); 
    assign layer_0[11344] = ~(in[788] ^ in[65]); 
    assign layer_0[11345] = ~in[998] | (in[998] & in[824]); 
    assign layer_0[11346] = in[504] & in[588]; 
    assign layer_0[11347] = ~in[652] | (in[754] & in[652]); 
    assign layer_0[11348] = ~(in[603] ^ in[668]); 
    assign layer_0[11349] = in[475] & ~in[922]; 
    assign layer_0[11350] = in[886] & in[872]; 
    assign layer_0[11351] = in[976] & ~in[859]; 
    assign layer_0[11352] = 1'b0; 
    assign layer_0[11353] = ~in[779] | (in[779] & in[783]); 
    assign layer_0[11354] = in[84] & in[950]; 
    assign layer_0[11355] = ~(in[299] ^ in[235]); 
    assign layer_0[11356] = ~(in[789] | in[18]); 
    assign layer_0[11357] = ~(in[744] ^ in[408]); 
    assign layer_0[11358] = in[776] ^ in[68]; 
    assign layer_0[11359] = in[600] & ~in[225]; 
    assign layer_0[11360] = in[845] & ~in[306]; 
    assign layer_0[11361] = in[604]; 
    assign layer_0[11362] = in[934] & ~in[802]; 
    assign layer_0[11363] = ~in[59]; 
    assign layer_0[11364] = in[876] ^ in[841]; 
    assign layer_0[11365] = ~in[124] | (in[124] & in[830]); 
    assign layer_0[11366] = in[102]; 
    assign layer_0[11367] = in[646]; 
    assign layer_0[11368] = ~(in[618] ^ in[597]); 
    assign layer_0[11369] = ~(in[93] & in[887]); 
    assign layer_0[11370] = in[12] & ~in[126]; 
    assign layer_0[11371] = ~in[906] | (in[906] & in[234]); 
    assign layer_0[11372] = in[410] & ~in[542]; 
    assign layer_0[11373] = in[244] | in[162]; 
    assign layer_0[11374] = in[20] | in[632]; 
    assign layer_0[11375] = ~(in[9] & in[711]); 
    assign layer_0[11376] = ~(in[550] & in[267]); 
    assign layer_0[11377] = ~in[857]; 
    assign layer_0[11378] = ~in[689]; 
    assign layer_0[11379] = ~(in[43] ^ in[854]); 
    assign layer_0[11380] = in[499] ^ in[954]; 
    assign layer_0[11381] = in[125] ^ in[11]; 
    assign layer_0[11382] = ~(in[549] ^ in[178]); 
    assign layer_0[11383] = in[821] & in[803]; 
    assign layer_0[11384] = in[932] & ~in[45]; 
    assign layer_0[11385] = ~(in[307] ^ in[589]); 
    assign layer_0[11386] = in[953] & in[826]; 
    assign layer_0[11387] = in[874] & ~in[793]; 
    assign layer_0[11388] = ~in[633] | (in[633] & in[192]); 
    assign layer_0[11389] = ~in[600] | (in[600] & in[763]); 
    assign layer_0[11390] = in[145] & ~in[132]; 
    assign layer_0[11391] = ~in[461]; 
    assign layer_0[11392] = in[428] & ~in[33]; 
    assign layer_0[11393] = in[713] | in[848]; 
    assign layer_0[11394] = in[157]; 
    assign layer_0[11395] = ~in[461]; 
    assign layer_0[11396] = ~(in[473] ^ in[598]); 
    assign layer_0[11397] = in[385] ^ in[595]; 
    assign layer_0[11398] = ~(in[339] & in[36]); 
    assign layer_0[11399] = in[499] ^ in[61]; 
    assign layer_0[11400] = in[1001] ^ in[93]; 
    assign layer_0[11401] = in[311]; 
    assign layer_0[11402] = in[666] ^ in[712]; 
    assign layer_0[11403] = ~(in[194] ^ in[983]); 
    assign layer_0[11404] = ~in[363]; 
    assign layer_0[11405] = ~(in[588] | in[955]); 
    assign layer_0[11406] = ~(in[437] & in[536]); 
    assign layer_0[11407] = in[445]; 
    assign layer_0[11408] = in[671] & in[955]; 
    assign layer_0[11409] = ~(in[974] ^ in[632]); 
    assign layer_0[11410] = ~(in[287] | in[627]); 
    assign layer_0[11411] = in[840]; 
    assign layer_0[11412] = ~(in[791] & in[665]); 
    assign layer_0[11413] = ~in[156]; 
    assign layer_0[11414] = in[554]; 
    assign layer_0[11415] = ~in[819]; 
    assign layer_0[11416] = ~in[140]; 
    assign layer_0[11417] = ~in[500] | (in[687] & in[500]); 
    assign layer_0[11418] = in[722] & in[709]; 
    assign layer_0[11419] = in[379]; 
    assign layer_0[11420] = in[1006] & ~in[35]; 
    assign layer_0[11421] = ~in[693]; 
    assign layer_0[11422] = in[757] | in[553]; 
    assign layer_0[11423] = ~in[538] | (in[538] & in[1015]); 
    assign layer_0[11424] = ~(in[930] & in[900]); 
    assign layer_0[11425] = ~in[471]; 
    assign layer_0[11426] = ~in[807] | (in[367] & in[807]); 
    assign layer_0[11427] = in[483] | in[654]; 
    assign layer_0[11428] = ~in[554] | (in[554] & in[889]); 
    assign layer_0[11429] = ~(in[533] & in[551]); 
    assign layer_0[11430] = ~(in[83] ^ in[62]); 
    assign layer_0[11431] = in[191] | in[259]; 
    assign layer_0[11432] = ~(in[747] ^ in[827]); 
    assign layer_0[11433] = in[694] ^ in[345]; 
    assign layer_0[11434] = ~in[613] | (in[613] & in[462]); 
    assign layer_0[11435] = ~(in[84] ^ in[442]); 
    assign layer_0[11436] = in[344]; 
    assign layer_0[11437] = in[640] ^ in[570]; 
    assign layer_0[11438] = ~(in[668] ^ in[915]); 
    assign layer_0[11439] = ~in[44]; 
    assign layer_0[11440] = ~in[126]; 
    assign layer_0[11441] = ~(in[931] & in[193]); 
    assign layer_0[11442] = in[553] | in[860]; 
    assign layer_0[11443] = ~(in[705] ^ in[177]); 
    assign layer_0[11444] = ~in[477] | (in[477] & in[759]); 
    assign layer_0[11445] = ~(in[632] ^ in[744]); 
    assign layer_0[11446] = ~(in[232] ^ in[45]); 
    assign layer_0[11447] = ~(in[146] & in[146]); 
    assign layer_0[11448] = ~(in[185] & in[632]); 
    assign layer_0[11449] = ~(in[118] ^ in[308]); 
    assign layer_0[11450] = ~in[586] | (in[586] & in[258]); 
    assign layer_0[11451] = ~(in[29] ^ in[635]); 
    assign layer_0[11452] = in[749] ^ in[659]; 
    assign layer_0[11453] = ~(in[597] & in[602]); 
    assign layer_0[11454] = in[614] | in[248]; 
    assign layer_0[11455] = in[787]; 
    assign layer_0[11456] = in[700]; 
    assign layer_0[11457] = ~(in[992] & in[650]); 
    assign layer_0[11458] = ~(in[614] ^ in[941]); 
    assign layer_0[11459] = ~in[766] | (in[233] & in[766]); 
    assign layer_0[11460] = in[843] ^ in[855]; 
    assign layer_0[11461] = in[470]; 
    assign layer_0[11462] = ~(in[706] & in[405]); 
    assign layer_0[11463] = in[937]; 
    assign layer_0[11464] = in[539] & in[10]; 
    assign layer_0[11465] = in[252] & in[296]; 
    assign layer_0[11466] = in[180] ^ in[225]; 
    assign layer_0[11467] = in[501] ^ in[108]; 
    assign layer_0[11468] = in[693] & in[589]; 
    assign layer_0[11469] = 1'b1; 
    assign layer_0[11470] = in[108]; 
    assign layer_0[11471] = in[308] ^ in[267]; 
    assign layer_0[11472] = in[675] | in[901]; 
    assign layer_0[11473] = ~(in[869] ^ in[583]); 
    assign layer_0[11474] = in[921] | in[854]; 
    assign layer_0[11475] = ~(in[886] & in[872]); 
    assign layer_0[11476] = 1'b1; 
    assign layer_0[11477] = in[548]; 
    assign layer_0[11478] = ~in[317]; 
    assign layer_0[11479] = ~in[981] | (in[981] & in[1001]); 
    assign layer_0[11480] = ~(in[699] ^ in[838]); 
    assign layer_0[11481] = ~(in[804] ^ in[595]); 
    assign layer_0[11482] = in[849]; 
    assign layer_0[11483] = in[448] | in[636]; 
    assign layer_0[11484] = ~in[553] | (in[542] & in[553]); 
    assign layer_0[11485] = in[290] ^ in[746]; 
    assign layer_0[11486] = in[974] | in[734]; 
    assign layer_0[11487] = ~(in[984] & in[550]); 
    assign layer_0[11488] = ~in[770] | (in[196] & in[770]); 
    assign layer_0[11489] = in[740] ^ in[249]; 
    assign layer_0[11490] = ~(in[918] & in[435]); 
    assign layer_0[11491] = in[79]; 
    assign layer_0[11492] = ~in[555] | (in[916] & in[555]); 
    assign layer_0[11493] = ~(in[806] ^ in[705]); 
    assign layer_0[11494] = ~(in[727] | in[956]); 
    assign layer_0[11495] = ~(in[91] ^ in[711]); 
    assign layer_0[11496] = ~(in[402] ^ in[794]); 
    assign layer_0[11497] = in[694] & in[311]; 
    assign layer_0[11498] = in[81] ^ in[925]; 
    assign layer_0[11499] = in[469]; 
    assign layer_0[11500] = ~(in[236] ^ in[211]); 
    assign layer_0[11501] = ~in[1014]; 
    assign layer_0[11502] = ~(in[518] | in[449]); 
    assign layer_0[11503] = ~(in[603] ^ in[698]); 
    assign layer_0[11504] = ~(in[856] ^ in[859]); 
    assign layer_0[11505] = in[893] ^ in[905]; 
    assign layer_0[11506] = in[219] & in[215]; 
    assign layer_0[11507] = in[719] & ~in[791]; 
    assign layer_0[11508] = ~in[697]; 
    assign layer_0[11509] = in[253] & in[26]; 
    assign layer_0[11510] = in[316] ^ in[11]; 
    assign layer_0[11511] = in[167] & ~in[607]; 
    assign layer_0[11512] = ~(in[582] ^ in[836]); 
    assign layer_0[11513] = ~(in[890] ^ in[970]); 
    assign layer_0[11514] = ~(in[605] | in[24]); 
    assign layer_0[11515] = in[824]; 
    assign layer_0[11516] = 1'b0; 
    assign layer_0[11517] = ~(in[484] ^ in[277]); 
    assign layer_0[11518] = in[155] & ~in[952]; 
    assign layer_0[11519] = 1'b1; 
    assign layer_0[11520] = in[692] ^ in[604]; 
    assign layer_0[11521] = in[659]; 
    assign layer_0[11522] = ~in[79]; 
    assign layer_0[11523] = in[461] ^ in[109]; 
    assign layer_0[11524] = ~in[130] | (in[910] & in[130]); 
    assign layer_0[11525] = ~(in[612] & in[598]); 
    assign layer_0[11526] = in[349] ^ in[504]; 
    assign layer_0[11527] = in[746] ^ in[1000]; 
    assign layer_0[11528] = in[642] | in[795]; 
    assign layer_0[11529] = in[572] ^ in[793]; 
    assign layer_0[11530] = in[472] & ~in[647]; 
    assign layer_0[11531] = in[693] & in[307]; 
    assign layer_0[11532] = in[379] & in[859]; 
    assign layer_0[11533] = in[1015] ^ in[434]; 
    assign layer_0[11534] = ~in[445]; 
    assign layer_0[11535] = ~(in[602] ^ in[947]); 
    assign layer_0[11536] = in[884] & ~in[873]; 
    assign layer_0[11537] = ~(in[393] & in[83]); 
    assign layer_0[11538] = ~(in[998] ^ in[411]); 
    assign layer_0[11539] = ~in[884] | (in[884] & in[184]); 
    assign layer_0[11540] = ~(in[230] ^ in[477]); 
    assign layer_0[11541] = in[901]; 
    assign layer_0[11542] = ~in[522]; 
    assign layer_0[11543] = ~(in[265] | in[78]); 
    assign layer_0[11544] = ~(in[39] ^ in[704]); 
    assign layer_0[11545] = in[821] | in[936]; 
    assign layer_0[11546] = ~(in[881] | in[1]); 
    assign layer_0[11547] = ~(in[853] ^ in[709]); 
    assign layer_0[11548] = in[853] & ~in[380]; 
    assign layer_0[11549] = ~in[397] | (in[397] & in[111]); 
    assign layer_0[11550] = ~(in[915] ^ in[701]); 
    assign layer_0[11551] = in[254] & ~in[283]; 
    assign layer_0[11552] = in[76] ^ in[36]; 
    assign layer_0[11553] = in[123] & in[179]; 
    assign layer_0[11554] = in[565] & ~in[787]; 
    assign layer_0[11555] = ~(in[7] ^ in[733]); 
    assign layer_0[11556] = ~(in[71] ^ in[315]); 
    assign layer_0[11557] = ~(in[898] ^ in[909]); 
    assign layer_0[11558] = ~in[666] | (in[666] & in[862]); 
    assign layer_0[11559] = ~(in[836] | in[603]); 
    assign layer_0[11560] = ~(in[569] & in[284]); 
    assign layer_0[11561] = in[1014] & ~in[80]; 
    assign layer_0[11562] = ~(in[759] | in[491]); 
    assign layer_0[11563] = 1'b0; 
    assign layer_0[11564] = in[437] ^ in[978]; 
    assign layer_0[11565] = ~(in[712] ^ in[574]); 
    assign layer_0[11566] = in[629] | in[32]; 
    assign layer_0[11567] = in[1020]; 
    assign layer_0[11568] = in[34] | in[361]; 
    assign layer_0[11569] = in[284]; 
    assign layer_0[11570] = in[427] & ~in[874]; 
    assign layer_0[11571] = ~in[458]; 
    assign layer_0[11572] = in[791] & ~in[253]; 
    assign layer_0[11573] = in[1012] ^ in[30]; 
    assign layer_0[11574] = in[672] ^ in[745]; 
    assign layer_0[11575] = ~in[604]; 
    assign layer_0[11576] = in[307] ^ in[992]; 
    assign layer_0[11577] = in[132] & ~in[921]; 
    assign layer_0[11578] = in[727] & ~in[104]; 
    assign layer_0[11579] = ~(in[636] ^ in[121]); 
    assign layer_0[11580] = in[62] | in[567]; 
    assign layer_0[11581] = in[749] ^ in[733]; 
    assign layer_0[11582] = ~(in[82] | in[532]); 
    assign layer_0[11583] = in[180] & in[488]; 
    assign layer_0[11584] = ~in[984] | (in[984] & in[959]); 
    assign layer_0[11585] = in[808] ^ in[736]; 
    assign layer_0[11586] = ~in[983] | (in[983] & in[522]); 
    assign layer_0[11587] = in[578] ^ in[763]; 
    assign layer_0[11588] = ~(in[909] | in[80]); 
    assign layer_0[11589] = in[764] ^ in[937]; 
    assign layer_0[11590] = in[468] ^ in[397]; 
    assign layer_0[11591] = in[997]; 
    assign layer_0[11592] = ~(in[197] ^ in[111]); 
    assign layer_0[11593] = ~in[655]; 
    assign layer_0[11594] = in[869] | in[948]; 
    assign layer_0[11595] = ~in[520] | (in[968] & in[520]); 
    assign layer_0[11596] = in[539] | in[640]; 
    assign layer_0[11597] = in[787]; 
    assign layer_0[11598] = ~(in[708] ^ in[868]); 
    assign layer_0[11599] = ~(in[979] | in[697]); 
    assign layer_0[11600] = ~(in[237] ^ in[635]); 
    assign layer_0[11601] = ~(in[531] ^ in[283]); 
    assign layer_0[11602] = in[1014]; 
    assign layer_0[11603] = in[184] & ~in[708]; 
    assign layer_0[11604] = in[979] ^ in[465]; 
    assign layer_0[11605] = ~(in[635] | in[724]); 
    assign layer_0[11606] = ~(in[616] ^ in[617]); 
    assign layer_0[11607] = in[910] & in[346]; 
    assign layer_0[11608] = in[602] ^ in[665]; 
    assign layer_0[11609] = in[746]; 
    assign layer_0[11610] = ~(in[625] ^ in[179]); 
    assign layer_0[11611] = ~in[875] | (in[875] & in[290]); 
    assign layer_0[11612] = 1'b1; 
    assign layer_0[11613] = in[74] ^ in[56]; 
    assign layer_0[11614] = ~(in[869] & in[565]); 
    assign layer_0[11615] = in[605]; 
    assign layer_0[11616] = ~in[911]; 
    assign layer_0[11617] = in[364] & in[60]; 
    assign layer_0[11618] = in[812] ^ in[861]; 
    assign layer_0[11619] = ~(in[79] ^ in[845]); 
    assign layer_0[11620] = in[105] & in[982]; 
    assign layer_0[11621] = ~(in[396] ^ in[853]); 
    assign layer_0[11622] = ~in[852]; 
    assign layer_0[11623] = in[550] & ~in[556]; 
    assign layer_0[11624] = ~(in[279] ^ in[177]); 
    assign layer_0[11625] = ~(in[523] ^ in[1001]); 
    assign layer_0[11626] = ~(in[663] ^ in[923]); 
    assign layer_0[11627] = in[412]; 
    assign layer_0[11628] = in[821] ^ in[822]; 
    assign layer_0[11629] = in[204] ^ in[114]; 
    assign layer_0[11630] = ~in[975] | (in[975] & in[869]); 
    assign layer_0[11631] = ~(in[558] ^ in[130]); 
    assign layer_0[11632] = ~(in[446] ^ in[374]); 
    assign layer_0[11633] = in[555] ^ in[94]; 
    assign layer_0[11634] = in[823] ^ in[691]; 
    assign layer_0[11635] = in[45]; 
    assign layer_0[11636] = in[582] & ~in[29]; 
    assign layer_0[11637] = ~(in[945] | in[370]); 
    assign layer_0[11638] = ~(in[39] ^ in[953]); 
    assign layer_0[11639] = ~(in[173] ^ in[354]); 
    assign layer_0[11640] = ~in[140] | (in[140] & in[700]); 
    assign layer_0[11641] = ~(in[948] ^ in[586]); 
    assign layer_0[11642] = in[40] & ~in[238]; 
    assign layer_0[11643] = ~in[791] | (in[471] & in[791]); 
    assign layer_0[11644] = in[0]; 
    assign layer_0[11645] = in[713] ^ in[878]; 
    assign layer_0[11646] = ~(in[383] ^ in[313]); 
    assign layer_0[11647] = in[921] & in[836]; 
    assign layer_0[11648] = in[660]; 
    assign layer_0[11649] = in[842]; 
    assign layer_0[11650] = ~(in[98] & in[884]); 
    assign layer_0[11651] = ~(in[605] ^ in[582]); 
    assign layer_0[11652] = ~(in[4] ^ in[500]); 
    assign layer_0[11653] = ~(in[1021] ^ in[334]); 
    assign layer_0[11654] = in[857] ^ in[858]; 
    assign layer_0[11655] = ~in[15]; 
    assign layer_0[11656] = ~(in[155] & in[604]); 
    assign layer_0[11657] = in[932] ^ in[128]; 
    assign layer_0[11658] = ~(in[554] ^ in[551]); 
    assign layer_0[11659] = ~(in[661] ^ in[29]); 
    assign layer_0[11660] = in[903] & ~in[833]; 
    assign layer_0[11661] = ~(in[613] & in[433]); 
    assign layer_0[11662] = in[475] & ~in[943]; 
    assign layer_0[11663] = ~(in[707] ^ in[238]); 
    assign layer_0[11664] = in[702]; 
    assign layer_0[11665] = ~in[190] | (in[190] & in[561]); 
    assign layer_0[11666] = in[711]; 
    assign layer_0[11667] = ~(in[650] & in[198]); 
    assign layer_0[11668] = in[25] | in[49]; 
    assign layer_0[11669] = ~(in[982] | in[517]); 
    assign layer_0[11670] = in[88] & ~in[744]; 
    assign layer_0[11671] = in[597] & ~in[1003]; 
    assign layer_0[11672] = in[182] ^ in[383]; 
    assign layer_0[11673] = ~(in[868] ^ in[412]); 
    assign layer_0[11674] = in[967] | in[657]; 
    assign layer_0[11675] = ~(in[953] | in[927]); 
    assign layer_0[11676] = ~in[673] | (in[673] & in[816]); 
    assign layer_0[11677] = ~in[726] | (in[927] & in[726]); 
    assign layer_0[11678] = in[60] & ~in[180]; 
    assign layer_0[11679] = in[174] ^ in[1016]; 
    assign layer_0[11680] = ~in[667] | (in[806] & in[667]); 
    assign layer_0[11681] = in[582] | in[719]; 
    assign layer_0[11682] = ~in[178] | (in[895] & in[178]); 
    assign layer_0[11683] = 1'b0; 
    assign layer_0[11684] = in[563] | in[290]; 
    assign layer_0[11685] = in[761] & ~in[415]; 
    assign layer_0[11686] = in[201] & ~in[221]; 
    assign layer_0[11687] = ~(in[345] & in[753]); 
    assign layer_0[11688] = in[98]; 
    assign layer_0[11689] = ~in[688]; 
    assign layer_0[11690] = in[588]; 
    assign layer_0[11691] = in[414] | in[449]; 
    assign layer_0[11692] = in[145] & ~in[580]; 
    assign layer_0[11693] = ~in[469] | (in[469] & in[433]); 
    assign layer_0[11694] = ~(in[358] ^ in[393]); 
    assign layer_0[11695] = in[870]; 
    assign layer_0[11696] = in[732] ^ in[940]; 
    assign layer_0[11697] = in[436] ^ in[952]; 
    assign layer_0[11698] = ~(in[403] ^ in[492]); 
    assign layer_0[11699] = in[308] & in[299]; 
    assign layer_0[11700] = in[196] ^ in[644]; 
    assign layer_0[11701] = ~in[566]; 
    assign layer_0[11702] = ~in[586] | (in[586] & in[355]); 
    assign layer_0[11703] = in[29] ^ in[241]; 
    assign layer_0[11704] = in[914]; 
    assign layer_0[11705] = ~(in[729] ^ in[587]); 
    assign layer_0[11706] = ~in[573]; 
    assign layer_0[11707] = in[229] ^ in[315]; 
    assign layer_0[11708] = in[808] | in[784]; 
    assign layer_0[11709] = in[209] & in[954]; 
    assign layer_0[11710] = ~in[648] | (in[648] & in[813]); 
    assign layer_0[11711] = ~(in[570] ^ in[318]); 
    assign layer_0[11712] = ~in[170] | (in[504] & in[170]); 
    assign layer_0[11713] = in[631] ^ in[498]; 
    assign layer_0[11714] = in[3] | in[937]; 
    assign layer_0[11715] = ~(in[522] & in[949]); 
    assign layer_0[11716] = in[899] | in[974]; 
    assign layer_0[11717] = in[656] ^ in[791]; 
    assign layer_0[11718] = in[729] ^ in[318]; 
    assign layer_0[11719] = in[1015] | in[619]; 
    assign layer_0[11720] = in[146] ^ in[862]; 
    assign layer_0[11721] = in[958] ^ in[920]; 
    assign layer_0[11722] = ~in[583] | (in[3] & in[583]); 
    assign layer_0[11723] = 1'b1; 
    assign layer_0[11724] = ~(in[855] & in[922]); 
    assign layer_0[11725] = ~(in[335] ^ in[871]); 
    assign layer_0[11726] = ~(in[965] ^ in[870]); 
    assign layer_0[11727] = ~in[967]; 
    assign layer_0[11728] = in[381] & in[706]; 
    assign layer_0[11729] = ~(in[608] ^ in[25]); 
    assign layer_0[11730] = ~in[226] | (in[226] & in[900]); 
    assign layer_0[11731] = in[987] | in[238]; 
    assign layer_0[11732] = in[47] & ~in[172]; 
    assign layer_0[11733] = ~(in[351] & in[677]); 
    assign layer_0[11734] = in[961] | in[49]; 
    assign layer_0[11735] = ~in[604]; 
    assign layer_0[11736] = in[910] ^ in[252]; 
    assign layer_0[11737] = ~(in[162] & in[677]); 
    assign layer_0[11738] = in[984] & ~in[835]; 
    assign layer_0[11739] = ~(in[953] & in[965]); 
    assign layer_0[11740] = in[507] | in[500]; 
    assign layer_0[11741] = in[223] ^ in[159]; 
    assign layer_0[11742] = ~(in[41] & in[386]); 
    assign layer_0[11743] = in[397] & ~in[644]; 
    assign layer_0[11744] = ~(in[480] | in[416]); 
    assign layer_0[11745] = in[81] ^ in[706]; 
    assign layer_0[11746] = ~in[116]; 
    assign layer_0[11747] = ~in[585]; 
    assign layer_0[11748] = in[696] & in[460]; 
    assign layer_0[11749] = in[435] & ~in[478]; 
    assign layer_0[11750] = ~(in[363] & in[632]); 
    assign layer_0[11751] = ~(in[222] & in[489]); 
    assign layer_0[11752] = in[58] ^ in[911]; 
    assign layer_0[11753] = ~in[195]; 
    assign layer_0[11754] = in[363] & in[596]; 
    assign layer_0[11755] = ~in[684] | (in[684] & in[498]); 
    assign layer_0[11756] = ~(in[208] & in[600]); 
    assign layer_0[11757] = in[521] & ~in[956]; 
    assign layer_0[11758] = 1'b0; 
    assign layer_0[11759] = in[207]; 
    assign layer_0[11760] = in[314] ^ in[733]; 
    assign layer_0[11761] = ~in[281] | (in[17] & in[281]); 
    assign layer_0[11762] = in[756] | in[317]; 
    assign layer_0[11763] = ~(in[709] & in[602]); 
    assign layer_0[11764] = in[689] ^ in[355]; 
    assign layer_0[11765] = ~(in[216] | in[95]); 
    assign layer_0[11766] = ~(in[570] ^ in[810]); 
    assign layer_0[11767] = in[220] ^ in[695]; 
    assign layer_0[11768] = in[261] ^ in[293]; 
    assign layer_0[11769] = ~(in[869] ^ in[981]); 
    assign layer_0[11770] = in[813] ^ in[956]; 
    assign layer_0[11771] = in[606] ^ in[145]; 
    assign layer_0[11772] = in[319] ^ in[702]; 
    assign layer_0[11773] = ~in[492] | (in[492] & in[461]); 
    assign layer_0[11774] = ~in[447]; 
    assign layer_0[11775] = in[198] & ~in[759]; 
    assign layer_0[11776] = ~(in[859] & in[56]); 
    assign layer_0[11777] = in[550] | in[445]; 
    assign layer_0[11778] = in[108] ^ in[756]; 
    assign layer_0[11779] = ~(in[819] | in[909]); 
    assign layer_0[11780] = in[823] ^ in[993]; 
    assign layer_0[11781] = in[228]; 
    assign layer_0[11782] = in[24] & in[737]; 
    assign layer_0[11783] = ~(in[794] ^ in[791]); 
    assign layer_0[11784] = in[954] ^ in[124]; 
    assign layer_0[11785] = in[926] & ~in[719]; 
    assign layer_0[11786] = in[607]; 
    assign layer_0[11787] = in[599]; 
    assign layer_0[11788] = in[823] ^ in[822]; 
    assign layer_0[11789] = ~(in[242] ^ in[347]); 
    assign layer_0[11790] = in[212] & ~in[941]; 
    assign layer_0[11791] = ~(in[242] & in[50]); 
    assign layer_0[11792] = ~(in[999] ^ in[790]); 
    assign layer_0[11793] = ~(in[489] | in[612]); 
    assign layer_0[11794] = ~(in[767] ^ in[20]); 
    assign layer_0[11795] = in[517] ^ in[401]; 
    assign layer_0[11796] = in[389] & ~in[931]; 
    assign layer_0[11797] = in[882]; 
    assign layer_0[11798] = 1'b0; 
    assign layer_0[11799] = in[428] ^ in[476]; 
    assign layer_0[11800] = in[900] | in[195]; 
    assign layer_0[11801] = in[677]; 
    assign layer_0[11802] = ~(in[914] ^ in[983]); 
    assign layer_0[11803] = ~in[392]; 
    assign layer_0[11804] = ~(in[268] ^ in[189]); 
    assign layer_0[11805] = ~(in[661] | in[234]); 
    assign layer_0[11806] = 1'b0; 
    assign layer_0[11807] = in[331] ^ in[965]; 
    assign layer_0[11808] = ~(in[301] | in[999]); 
    assign layer_0[11809] = in[218] & ~in[332]; 
    assign layer_0[11810] = ~in[340]; 
    assign layer_0[11811] = in[537] ^ in[885]; 
    assign layer_0[11812] = in[552] ^ in[553]; 
    assign layer_0[11813] = ~(in[513] ^ in[100]); 
    assign layer_0[11814] = in[551] & ~in[261]; 
    assign layer_0[11815] = 1'b0; 
    assign layer_0[11816] = ~in[710] | (in[710] & in[870]); 
    assign layer_0[11817] = ~(in[886] ^ in[853]); 
    assign layer_0[11818] = ~in[927]; 
    assign layer_0[11819] = in[581]; 
    assign layer_0[11820] = ~(in[67] | in[564]); 
    assign layer_0[11821] = ~(in[1000] ^ in[603]); 
    assign layer_0[11822] = ~(in[568] ^ in[28]); 
    assign layer_0[11823] = in[333] & ~in[998]; 
    assign layer_0[11824] = ~in[427] | (in[734] & in[427]); 
    assign layer_0[11825] = ~(in[120] ^ in[572]); 
    assign layer_0[11826] = in[822] & ~in[300]; 
    assign layer_0[11827] = in[871] ^ in[605]; 
    assign layer_0[11828] = ~(in[641] ^ in[794]); 
    assign layer_0[11829] = ~(in[886] ^ in[871]); 
    assign layer_0[11830] = ~in[171]; 
    assign layer_0[11831] = in[933] | in[921]; 
    assign layer_0[11832] = ~(in[792] | in[809]); 
    assign layer_0[11833] = ~(in[661] | in[1017]); 
    assign layer_0[11834] = ~(in[992] ^ in[643]); 
    assign layer_0[11835] = ~in[872]; 
    assign layer_0[11836] = ~in[11]; 
    assign layer_0[11837] = ~in[404] | (in[404] & in[767]); 
    assign layer_0[11838] = ~in[426] | (in[426] & in[867]); 
    assign layer_0[11839] = ~(in[144] ^ in[868]); 
    assign layer_0[11840] = ~in[55] | (in[55] & in[271]); 
    assign layer_0[11841] = ~in[871]; 
    assign layer_0[11842] = in[942] | in[234]; 
    assign layer_0[11843] = in[931] | in[536]; 
    assign layer_0[11844] = in[980] | in[110]; 
    assign layer_0[11845] = ~(in[495] & in[31]); 
    assign layer_0[11846] = 1'b0; 
    assign layer_0[11847] = in[168]; 
    assign layer_0[11848] = ~in[908] | (in[545] & in[908]); 
    assign layer_0[11849] = in[829]; 
    assign layer_0[11850] = ~(in[627] ^ in[929]); 
    assign layer_0[11851] = ~in[2]; 
    assign layer_0[11852] = ~in[396] | (in[206] & in[396]); 
    assign layer_0[11853] = in[298] & ~in[492]; 
    assign layer_0[11854] = in[856] & ~in[591]; 
    assign layer_0[11855] = in[310]; 
    assign layer_0[11856] = in[160] & ~in[774]; 
    assign layer_0[11857] = in[403] & ~in[706]; 
    assign layer_0[11858] = ~in[339] | (in[339] & in[19]); 
    assign layer_0[11859] = in[929] | in[930]; 
    assign layer_0[11860] = in[424] & in[364]; 
    assign layer_0[11861] = in[387] ^ in[321]; 
    assign layer_0[11862] = ~(in[523] ^ in[119]); 
    assign layer_0[11863] = ~in[602] | (in[811] & in[602]); 
    assign layer_0[11864] = in[78] | in[977]; 
    assign layer_0[11865] = in[665] ^ in[664]; 
    assign layer_0[11866] = in[616] & in[442]; 
    assign layer_0[11867] = in[324] ^ in[654]; 
    assign layer_0[11868] = in[252] & in[44]; 
    assign layer_0[11869] = ~(in[835] ^ in[261]); 
    assign layer_0[11870] = ~(in[268] ^ in[683]); 
    assign layer_0[11871] = ~in[329] | (in[329] & in[563]); 
    assign layer_0[11872] = in[746] & ~in[314]; 
    assign layer_0[11873] = ~(in[241] ^ in[252]); 
    assign layer_0[11874] = ~in[824]; 
    assign layer_0[11875] = ~in[86] | (in[568] & in[86]); 
    assign layer_0[11876] = in[292] ^ in[347]; 
    assign layer_0[11877] = ~(in[552] ^ in[824]); 
    assign layer_0[11878] = in[866] ^ in[961]; 
    assign layer_0[11879] = in[113] ^ in[874]; 
    assign layer_0[11880] = in[792] ^ in[981]; 
    assign layer_0[11881] = in[715] ^ in[844]; 
    assign layer_0[11882] = ~(in[725] & in[248]); 
    assign layer_0[11883] = ~(in[213] ^ in[1016]); 
    assign layer_0[11884] = ~(in[947] | in[614]); 
    assign layer_0[11885] = ~in[488]; 
    assign layer_0[11886] = ~in[910]; 
    assign layer_0[11887] = in[870] ^ in[927]; 
    assign layer_0[11888] = 1'b1; 
    assign layer_0[11889] = in[824] | in[635]; 
    assign layer_0[11890] = in[290] & ~in[779]; 
    assign layer_0[11891] = ~(in[882] ^ in[1017]); 
    assign layer_0[11892] = in[908] ^ in[574]; 
    assign layer_0[11893] = in[129] ^ in[261]; 
    assign layer_0[11894] = in[943] & ~in[911]; 
    assign layer_0[11895] = in[140] & in[520]; 
    assign layer_0[11896] = ~in[932] | (in[61] & in[932]); 
    assign layer_0[11897] = in[540] | in[522]; 
    assign layer_0[11898] = ~in[317] | (in[317] & in[607]); 
    assign layer_0[11899] = ~(in[133] & in[837]); 
    assign layer_0[11900] = ~(in[888] ^ in[965]); 
    assign layer_0[11901] = ~(in[666] ^ in[918]); 
    assign layer_0[11902] = in[1017] & ~in[1015]; 
    assign layer_0[11903] = ~(in[733] | in[1021]); 
    assign layer_0[11904] = ~(in[635] ^ in[804]); 
    assign layer_0[11905] = in[591] ^ in[628]; 
    assign layer_0[11906] = in[563] & ~in[499]; 
    assign layer_0[11907] = ~in[276] | (in[222] & in[276]); 
    assign layer_0[11908] = ~in[22] | (in[22] & in[463]); 
    assign layer_0[11909] = in[326]; 
    assign layer_0[11910] = in[555] & ~in[522]; 
    assign layer_0[11911] = in[362] & in[1023]; 
    assign layer_0[11912] = ~in[602] | (in[602] & in[980]); 
    assign layer_0[11913] = ~in[301] | (in[516] & in[301]); 
    assign layer_0[11914] = ~(in[676] & in[892]); 
    assign layer_0[11915] = in[316] & in[947]; 
    assign layer_0[11916] = ~in[460] | (in[460] & in[33]); 
    assign layer_0[11917] = ~in[982] | (in[982] & in[354]); 
    assign layer_0[11918] = ~in[267]; 
    assign layer_0[11919] = ~in[98] | (in[98] & in[793]); 
    assign layer_0[11920] = ~(in[125] & in[905]); 
    assign layer_0[11921] = ~(in[477] ^ in[99]); 
    assign layer_0[11922] = in[296] ^ in[5]; 
    assign layer_0[11923] = in[898] ^ in[309]; 
    assign layer_0[11924] = in[247] ^ in[725]; 
    assign layer_0[11925] = in[997] ^ in[614]; 
    assign layer_0[11926] = ~(in[551] ^ in[571]); 
    assign layer_0[11927] = ~in[283]; 
    assign layer_0[11928] = ~(in[679] & in[967]); 
    assign layer_0[11929] = ~(in[757] ^ in[236]); 
    assign layer_0[11930] = ~(in[689] ^ in[479]); 
    assign layer_0[11931] = in[730] ^ in[234]; 
    assign layer_0[11932] = in[84] ^ in[97]; 
    assign layer_0[11933] = ~(in[532] | in[195]); 
    assign layer_0[11934] = in[888] ^ in[870]; 
    assign layer_0[11935] = in[856] ^ in[934]; 
    assign layer_0[11936] = in[852] & in[164]; 
    assign layer_0[11937] = in[565] & ~in[317]; 
    assign layer_0[11938] = in[308] & in[690]; 
    assign layer_0[11939] = in[647] ^ in[711]; 
    assign layer_0[11940] = in[226] ^ in[570]; 
    assign layer_0[11941] = in[66] & ~in[801]; 
    assign layer_0[11942] = in[939] & in[98]; 
    assign layer_0[11943] = ~in[339]; 
    assign layer_0[11944] = in[229] & ~in[147]; 
    assign layer_0[11945] = in[591] ^ in[478]; 
    assign layer_0[11946] = in[571] ^ in[523]; 
    assign layer_0[11947] = in[952] ^ in[934]; 
    assign layer_0[11948] = in[969] ^ in[571]; 
    assign layer_0[11949] = in[262]; 
    assign layer_0[11950] = in[695] & ~in[604]; 
    assign layer_0[11951] = ~(in[907] ^ in[242]); 
    assign layer_0[11952] = ~(in[668] ^ in[602]); 
    assign layer_0[11953] = in[885]; 
    assign layer_0[11954] = ~(in[794] ^ in[851]); 
    assign layer_0[11955] = ~(in[694] | in[851]); 
    assign layer_0[11956] = ~in[569] | (in[780] & in[569]); 
    assign layer_0[11957] = ~in[707]; 
    assign layer_0[11958] = in[272] & in[135]; 
    assign layer_0[11959] = in[692] ^ in[252]; 
    assign layer_0[11960] = in[429]; 
    assign layer_0[11961] = in[695] & ~in[258]; 
    assign layer_0[11962] = in[830] | in[286]; 
    assign layer_0[11963] = ~in[20] | (in[20] & in[780]); 
    assign layer_0[11964] = in[178] & in[920]; 
    assign layer_0[11965] = ~in[473] | (in[473] & in[540]); 
    assign layer_0[11966] = in[183]; 
    assign layer_0[11967] = ~in[603] | (in[603] & in[508]); 
    assign layer_0[11968] = ~in[253] | (in[253] & in[183]); 
    assign layer_0[11969] = in[423] & ~in[389]; 
    assign layer_0[11970] = in[457]; 
    assign layer_0[11971] = ~(in[599] | in[80]); 
    assign layer_0[11972] = in[266] ^ in[264]; 
    assign layer_0[11973] = ~(in[317] ^ in[278]); 
    assign layer_0[11974] = in[708]; 
    assign layer_0[11975] = in[654] & in[633]; 
    assign layer_0[11976] = ~(in[704] | in[829]); 
    assign layer_0[11977] = in[722] ^ in[673]; 
    assign layer_0[11978] = in[489] ^ in[724]; 
    assign layer_0[11979] = in[1020] & ~in[36]; 
    assign layer_0[11980] = in[492] | in[989]; 
    assign layer_0[11981] = ~(in[948] ^ in[451]); 
    assign layer_0[11982] = in[807]; 
    assign layer_0[11983] = ~in[723] | (in[277] & in[723]); 
    assign layer_0[11984] = in[504] ^ in[370]; 
    assign layer_0[11985] = ~(in[294] | in[165]); 
    assign layer_0[11986] = in[507] ^ in[504]; 
    assign layer_0[11987] = ~(in[775] & in[548]); 
    assign layer_0[11988] = in[568] ^ in[579]; 
    assign layer_0[11989] = in[950]; 
    assign layer_0[11990] = ~in[7] | (in[466] & in[7]); 
    assign layer_0[11991] = in[984] ^ in[579]; 
    assign layer_0[11992] = in[264] ^ in[600]; 
    assign layer_0[11993] = ~(in[65] ^ in[138]); 
    assign layer_0[11994] = in[888] & ~in[237]; 
    assign layer_0[11995] = ~in[746] | (in[746] & in[731]); 
    assign layer_0[11996] = ~in[417] | (in[417] & in[1001]); 
    assign layer_0[11997] = ~(in[203] ^ in[224]); 
    assign layer_0[11998] = in[101] & in[65]; 
    assign layer_0[11999] = ~in[266]; 
    // Layer 1 ============================================================
    assign out[0] = ~(layer_0[9521] ^ layer_0[1370]); 
    assign out[1] = layer_0[7130] ^ layer_0[10899]; 
    assign out[2] = ~layer_0[1815]; 
    assign out[3] = ~layer_0[5560]; 
    assign out[4] = ~layer_0[5200] | (layer_0[6076] & layer_0[5200]); 
    assign out[5] = layer_0[10541] ^ layer_0[1826]; 
    assign out[6] = ~layer_0[10775] | (layer_0[2387] & layer_0[10775]); 
    assign out[7] = layer_0[1225] ^ layer_0[2055]; 
    assign out[8] = ~(layer_0[6538] | layer_0[10178]); 
    assign out[9] = layer_0[2956] ^ layer_0[6453]; 
    assign out[10] = layer_0[6572] ^ layer_0[5538]; 
    assign out[11] = layer_0[3208]; 
    assign out[12] = layer_0[1263] & layer_0[5354]; 
    assign out[13] = layer_0[10080]; 
    assign out[14] = ~layer_0[10184] | (layer_0[10184] & layer_0[11314]); 
    assign out[15] = layer_0[9901] | layer_0[7812]; 
    assign out[16] = ~(layer_0[9163] ^ layer_0[6270]); 
    assign out[17] = ~(layer_0[3061] ^ layer_0[3084]); 
    assign out[18] = ~(layer_0[2194] ^ layer_0[10871]); 
    assign out[19] = ~(layer_0[1342] ^ layer_0[6301]); 
    assign out[20] = layer_0[7467] & ~layer_0[2081]; 
    assign out[21] = layer_0[3558] ^ layer_0[8357]; 
    assign out[22] = ~(layer_0[3286] ^ layer_0[4783]); 
    assign out[23] = layer_0[6824] ^ layer_0[7418]; 
    assign out[24] = layer_0[6584] & layer_0[11556]; 
    assign out[25] = ~(layer_0[11998] ^ layer_0[4325]); 
    assign out[26] = ~(layer_0[4350] ^ layer_0[280]); 
    assign out[27] = ~(layer_0[7737] ^ layer_0[7144]); 
    assign out[28] = ~layer_0[8486]; 
    assign out[29] = layer_0[5722] ^ layer_0[8729]; 
    assign out[30] = ~(layer_0[5064] ^ layer_0[7372]); 
    assign out[31] = layer_0[1049]; 
    assign out[32] = layer_0[610] & ~layer_0[9593]; 
    assign out[33] = layer_0[5079] & ~layer_0[7022]; 
    assign out[34] = ~(layer_0[9905] ^ layer_0[6775]); 
    assign out[35] = layer_0[1108]; 
    assign out[36] = ~(layer_0[10436] ^ layer_0[3035]); 
    assign out[37] = layer_0[2348] ^ layer_0[10410]; 
    assign out[38] = ~layer_0[3227]; 
    assign out[39] = ~(layer_0[4173] ^ layer_0[1328]); 
    assign out[40] = layer_0[3693] & layer_0[2513]; 
    assign out[41] = ~(layer_0[11328] ^ layer_0[11139]); 
    assign out[42] = layer_0[8852] ^ layer_0[9766]; 
    assign out[43] = layer_0[5239] & layer_0[11073]; 
    assign out[44] = layer_0[9819] & ~layer_0[10485]; 
    assign out[45] = layer_0[8039]; 
    assign out[46] = ~(layer_0[7492] ^ layer_0[4749]); 
    assign out[47] = ~(layer_0[5036] ^ layer_0[6968]); 
    assign out[48] = layer_0[10952] ^ layer_0[116]; 
    assign out[49] = layer_0[4053] ^ layer_0[10357]; 
    assign out[50] = layer_0[6555] & ~layer_0[3978]; 
    assign out[51] = layer_0[6445] ^ layer_0[11178]; 
    assign out[52] = ~(layer_0[2773] ^ layer_0[4930]); 
    assign out[53] = layer_0[6873] ^ layer_0[10733]; 
    assign out[54] = ~(layer_0[3779] | layer_0[10040]); 
    assign out[55] = layer_0[8251] ^ layer_0[4603]; 
    assign out[56] = layer_0[3927] ^ layer_0[4475]; 
    assign out[57] = layer_0[1166] ^ layer_0[8898]; 
    assign out[58] = ~layer_0[1446]; 
    assign out[59] = ~(layer_0[10768] ^ layer_0[3236]); 
    assign out[60] = ~(layer_0[9401] ^ layer_0[6006]); 
    assign out[61] = ~layer_0[1314]; 
    assign out[62] = layer_0[9069] | layer_0[10255]; 
    assign out[63] = ~(layer_0[9348] & layer_0[3340]); 
    assign out[64] = layer_0[7383]; 
    assign out[65] = ~(layer_0[7212] ^ layer_0[2938]); 
    assign out[66] = layer_0[3419] ^ layer_0[8360]; 
    assign out[67] = layer_0[5143] ^ layer_0[10672]; 
    assign out[68] = ~(layer_0[10499] & layer_0[9266]); 
    assign out[69] = ~layer_0[2759] | (layer_0[2759] & layer_0[4658]); 
    assign out[70] = layer_0[1322] ^ layer_0[1550]; 
    assign out[71] = layer_0[8749] ^ layer_0[6201]; 
    assign out[72] = ~layer_0[9046]; 
    assign out[73] = layer_0[3209] ^ layer_0[4682]; 
    assign out[74] = ~(layer_0[2566] ^ layer_0[3079]); 
    assign out[75] = ~layer_0[4975]; 
    assign out[76] = ~(layer_0[11520] ^ layer_0[5241]); 
    assign out[77] = ~layer_0[10041] | (layer_0[10041] & layer_0[9638]); 
    assign out[78] = ~layer_0[2345]; 
    assign out[79] = layer_0[5743] ^ layer_0[7489]; 
    assign out[80] = layer_0[2619] ^ layer_0[3135]; 
    assign out[81] = layer_0[7177]; 
    assign out[82] = layer_0[4155] ^ layer_0[5715]; 
    assign out[83] = ~layer_0[11936] | (layer_0[415] & layer_0[11936]); 
    assign out[84] = layer_0[6906] ^ layer_0[5656]; 
    assign out[85] = layer_0[7549] | layer_0[6361]; 
    assign out[86] = layer_0[711] ^ layer_0[11861]; 
    assign out[87] = ~layer_0[8824]; 
    assign out[88] = layer_0[3163] ^ layer_0[8408]; 
    assign out[89] = ~(layer_0[10952] ^ layer_0[1999]); 
    assign out[90] = ~(layer_0[10385] ^ layer_0[1222]); 
    assign out[91] = ~(layer_0[2874] ^ layer_0[8211]); 
    assign out[92] = layer_0[480]; 
    assign out[93] = ~(layer_0[4978] ^ layer_0[4928]); 
    assign out[94] = layer_0[4935]; 
    assign out[95] = ~(layer_0[6875] & layer_0[6990]); 
    assign out[96] = ~(layer_0[6186] ^ layer_0[3256]); 
    assign out[97] = layer_0[2440] ^ layer_0[6510]; 
    assign out[98] = layer_0[6732] | layer_0[2960]; 
    assign out[99] = ~layer_0[7609]; 
    assign out[100] = ~(layer_0[8476] ^ layer_0[3293]); 
    assign out[101] = ~(layer_0[5505] ^ layer_0[6997]); 
    assign out[102] = layer_0[3594] & ~layer_0[11578]; 
    assign out[103] = layer_0[11600]; 
    assign out[104] = layer_0[6599] ^ layer_0[5914]; 
    assign out[105] = ~(layer_0[2104] ^ layer_0[11450]); 
    assign out[106] = ~layer_0[4424]; 
    assign out[107] = ~(layer_0[9374] ^ layer_0[7921]); 
    assign out[108] = layer_0[4417] ^ layer_0[9847]; 
    assign out[109] = layer_0[3954] ^ layer_0[5461]; 
    assign out[110] = layer_0[8387] ^ layer_0[11518]; 
    assign out[111] = layer_0[6111] ^ layer_0[9464]; 
    assign out[112] = ~(layer_0[410] ^ layer_0[5429]); 
    assign out[113] = ~(layer_0[7919] ^ layer_0[3119]); 
    assign out[114] = ~(layer_0[1769] ^ layer_0[11220]); 
    assign out[115] = layer_0[9789] & ~layer_0[7159]; 
    assign out[116] = layer_0[10187] ^ layer_0[1584]; 
    assign out[117] = ~(layer_0[5325] ^ layer_0[6652]); 
    assign out[118] = ~(layer_0[9217] & layer_0[6315]); 
    assign out[119] = ~(layer_0[4758] ^ layer_0[5346]); 
    assign out[120] = layer_0[3755] ^ layer_0[1383]; 
    assign out[121] = layer_0[5824] | layer_0[10484]; 
    assign out[122] = layer_0[10171] ^ layer_0[11878]; 
    assign out[123] = ~layer_0[3582] | (layer_0[3582] & layer_0[6199]); 
    assign out[124] = ~(layer_0[2892] ^ layer_0[2154]); 
    assign out[125] = ~layer_0[7805] | (layer_0[11554] & layer_0[7805]); 
    assign out[126] = layer_0[11766] ^ layer_0[8348]; 
    assign out[127] = layer_0[7042] & layer_0[11790]; 
    assign out[128] = ~(layer_0[928] ^ layer_0[6668]); 
    assign out[129] = layer_0[9662] ^ layer_0[11330]; 
    assign out[130] = layer_0[7130] ^ layer_0[722]; 
    assign out[131] = layer_0[11693] ^ layer_0[185]; 
    assign out[132] = layer_0[4671]; 
    assign out[133] = layer_0[2953] & ~layer_0[5164]; 
    assign out[134] = layer_0[11995]; 
    assign out[135] = ~(layer_0[6335] ^ layer_0[3916]); 
    assign out[136] = layer_0[8595] ^ layer_0[8949]; 
    assign out[137] = ~layer_0[1060]; 
    assign out[138] = layer_0[7033]; 
    assign out[139] = layer_0[9437] ^ layer_0[2842]; 
    assign out[140] = layer_0[5434] ^ layer_0[10958]; 
    assign out[141] = ~(layer_0[4961] ^ layer_0[5566]); 
    assign out[142] = ~layer_0[8529] | (layer_0[2476] & layer_0[8529]); 
    assign out[143] = layer_0[7839] | layer_0[9403]; 
    assign out[144] = ~(layer_0[7416] ^ layer_0[7111]); 
    assign out[145] = layer_0[10620] & layer_0[2646]; 
    assign out[146] = layer_0[4980] ^ layer_0[8174]; 
    assign out[147] = 1'b0; 
    assign out[148] = layer_0[588] & layer_0[684]; 
    assign out[149] = layer_0[1694]; 
    assign out[150] = layer_0[2189] ^ layer_0[2154]; 
    assign out[151] = ~(layer_0[5709] ^ layer_0[6513]); 
    assign out[152] = layer_0[11224]; 
    assign out[153] = layer_0[1502]; 
    assign out[154] = layer_0[5667] & ~layer_0[1112]; 
    assign out[155] = layer_0[6176] ^ layer_0[6423]; 
    assign out[156] = layer_0[2626] ^ layer_0[4955]; 
    assign out[157] = layer_0[5098] & ~layer_0[6771]; 
    assign out[158] = ~(layer_0[6279] ^ layer_0[5806]); 
    assign out[159] = layer_0[1998] & layer_0[9485]; 
    assign out[160] = layer_0[7824] ^ layer_0[2182]; 
    assign out[161] = layer_0[1494] ^ layer_0[3632]; 
    assign out[162] = ~layer_0[9586]; 
    assign out[163] = layer_0[10686]; 
    assign out[164] = ~(layer_0[6288] ^ layer_0[10972]); 
    assign out[165] = layer_0[10426] ^ layer_0[2268]; 
    assign out[166] = ~(layer_0[5246] & layer_0[7633]); 
    assign out[167] = ~layer_0[5343]; 
    assign out[168] = ~(layer_0[3893] ^ layer_0[2299]); 
    assign out[169] = layer_0[1387] ^ layer_0[10948]; 
    assign out[170] = layer_0[5417] & ~layer_0[5371]; 
    assign out[171] = ~(layer_0[11664] ^ layer_0[4936]); 
    assign out[172] = ~layer_0[4165]; 
    assign out[173] = layer_0[2985]; 
    assign out[174] = ~(layer_0[4618] & layer_0[2876]); 
    assign out[175] = ~(layer_0[2141] ^ layer_0[1753]); 
    assign out[176] = layer_0[207] ^ layer_0[795]; 
    assign out[177] = layer_0[10151] | layer_0[8187]; 
    assign out[178] = ~(layer_0[1315] ^ layer_0[11728]); 
    assign out[179] = ~(layer_0[2602] ^ layer_0[1564]); 
    assign out[180] = layer_0[9313] ^ layer_0[10373]; 
    assign out[181] = ~(layer_0[10104] ^ layer_0[8578]); 
    assign out[182] = ~(layer_0[10923] ^ layer_0[3382]); 
    assign out[183] = ~(layer_0[306] ^ layer_0[9835]); 
    assign out[184] = ~(layer_0[9552] ^ layer_0[4328]); 
    assign out[185] = layer_0[5594] & layer_0[7036]; 
    assign out[186] = layer_0[11807] ^ layer_0[774]; 
    assign out[187] = ~(layer_0[2530] | layer_0[5519]); 
    assign out[188] = layer_0[3474] ^ layer_0[5178]; 
    assign out[189] = layer_0[5359] & ~layer_0[5817]; 
    assign out[190] = ~(layer_0[4467] ^ layer_0[6408]); 
    assign out[191] = ~(layer_0[3587] ^ layer_0[5287]); 
    assign out[192] = layer_0[11849]; 
    assign out[193] = ~(layer_0[8746] ^ layer_0[4491]); 
    assign out[194] = ~(layer_0[11703] ^ layer_0[4866]); 
    assign out[195] = layer_0[7368] & ~layer_0[4545]; 
    assign out[196] = ~(layer_0[7108] ^ layer_0[4334]); 
    assign out[197] = ~(layer_0[6797] & layer_0[10683]); 
    assign out[198] = layer_0[1158]; 
    assign out[199] = ~(layer_0[11668] ^ layer_0[1178]); 
    assign out[200] = ~(layer_0[11895] ^ layer_0[6586]); 
    assign out[201] = layer_0[5034] ^ layer_0[9557]; 
    assign out[202] = ~(layer_0[4960] | layer_0[11788]); 
    assign out[203] = ~(layer_0[11585] ^ layer_0[7549]); 
    assign out[204] = ~(layer_0[9022] ^ layer_0[8834]); 
    assign out[205] = ~(layer_0[6066] ^ layer_0[4515]); 
    assign out[206] = layer_0[4587] & ~layer_0[1668]; 
    assign out[207] = ~(layer_0[9280] ^ layer_0[1029]); 
    assign out[208] = ~(layer_0[3168] ^ layer_0[11841]); 
    assign out[209] = layer_0[11874]; 
    assign out[210] = ~(layer_0[6164] ^ layer_0[4769]); 
    assign out[211] = ~(layer_0[4650] ^ layer_0[8378]); 
    assign out[212] = layer_0[6483] & layer_0[9399]; 
    assign out[213] = layer_0[825] ^ layer_0[11340]; 
    assign out[214] = ~layer_0[5893]; 
    assign out[215] = layer_0[3620] ^ layer_0[5831]; 
    assign out[216] = layer_0[3035] ^ layer_0[7550]; 
    assign out[217] = layer_0[5305]; 
    assign out[218] = ~layer_0[1627]; 
    assign out[219] = layer_0[1458] ^ layer_0[1579]; 
    assign out[220] = ~(layer_0[8867] & layer_0[881]); 
    assign out[221] = ~(layer_0[1114] ^ layer_0[1409]); 
    assign out[222] = ~(layer_0[9678] & layer_0[7912]); 
    assign out[223] = layer_0[10152] ^ layer_0[7533]; 
    assign out[224] = layer_0[5649] ^ layer_0[9361]; 
    assign out[225] = ~layer_0[7601]; 
    assign out[226] = ~layer_0[804]; 
    assign out[227] = layer_0[6405] & layer_0[130]; 
    assign out[228] = ~layer_0[5414]; 
    assign out[229] = layer_0[6531] ^ layer_0[8329]; 
    assign out[230] = ~(layer_0[3131] ^ layer_0[10925]); 
    assign out[231] = ~(layer_0[5622] ^ layer_0[8684]); 
    assign out[232] = ~(layer_0[9412] ^ layer_0[3984]); 
    assign out[233] = ~(layer_0[3025] ^ layer_0[5666]); 
    assign out[234] = layer_0[9971] & ~layer_0[10613]; 
    assign out[235] = layer_0[1943] & ~layer_0[7806]; 
    assign out[236] = ~(layer_0[6964] ^ layer_0[8088]); 
    assign out[237] = ~(layer_0[8173] ^ layer_0[6720]); 
    assign out[238] = layer_0[8736] ^ layer_0[3313]; 
    assign out[239] = layer_0[11829]; 
    assign out[240] = layer_0[9094] & layer_0[758]; 
    assign out[241] = layer_0[7626] ^ layer_0[5561]; 
    assign out[242] = layer_0[5855]; 
    assign out[243] = ~(layer_0[8396] ^ layer_0[6758]); 
    assign out[244] = ~(layer_0[4828] ^ layer_0[9723]); 
    assign out[245] = layer_0[2294] | layer_0[4555]; 
    assign out[246] = layer_0[3245] & ~layer_0[87]; 
    assign out[247] = ~(layer_0[8056] ^ layer_0[3714]); 
    assign out[248] = layer_0[5540]; 
    assign out[249] = layer_0[7718] ^ layer_0[5948]; 
    assign out[250] = ~layer_0[11436] | (layer_0[11436] & layer_0[1237]); 
    assign out[251] = layer_0[708] ^ layer_0[285]; 
    assign out[252] = layer_0[9422] ^ layer_0[8438]; 
    assign out[253] = ~(layer_0[10133] ^ layer_0[6811]); 
    assign out[254] = layer_0[2674] ^ layer_0[11470]; 
    assign out[255] = layer_0[591]; 
    assign out[256] = ~(layer_0[6698] ^ layer_0[1242]); 
    assign out[257] = ~(layer_0[8718] ^ layer_0[10872]); 
    assign out[258] = layer_0[10955] & ~layer_0[9607]; 
    assign out[259] = layer_0[1504] ^ layer_0[9483]; 
    assign out[260] = layer_0[7240] ^ layer_0[607]; 
    assign out[261] = ~layer_0[7655]; 
    assign out[262] = layer_0[5890] ^ layer_0[8794]; 
    assign out[263] = layer_0[5113] & layer_0[11203]; 
    assign out[264] = layer_0[3460] ^ layer_0[7621]; 
    assign out[265] = layer_0[10239] & ~layer_0[11432]; 
    assign out[266] = layer_0[8315] & ~layer_0[598]; 
    assign out[267] = layer_0[4521] & layer_0[2788]; 
    assign out[268] = ~(layer_0[7553] ^ layer_0[1244]); 
    assign out[269] = ~(layer_0[2957] ^ layer_0[8398]); 
    assign out[270] = layer_0[1211] ^ layer_0[2500]; 
    assign out[271] = ~(layer_0[8275] ^ layer_0[2504]); 
    assign out[272] = layer_0[4024] ^ layer_0[11038]; 
    assign out[273] = layer_0[7368] ^ layer_0[9990]; 
    assign out[274] = layer_0[8797] | layer_0[2440]; 
    assign out[275] = ~(layer_0[709] ^ layer_0[6230]); 
    assign out[276] = ~(layer_0[10627] ^ layer_0[3866]); 
    assign out[277] = ~(layer_0[4380] ^ layer_0[10267]); 
    assign out[278] = layer_0[903] ^ layer_0[9605]; 
    assign out[279] = ~layer_0[11205]; 
    assign out[280] = layer_0[10511] ^ layer_0[11386]; 
    assign out[281] = ~(layer_0[2778] ^ layer_0[780]); 
    assign out[282] = ~(layer_0[4549] ^ layer_0[5653]); 
    assign out[283] = layer_0[11914] & ~layer_0[7890]; 
    assign out[284] = ~(layer_0[9126] ^ layer_0[8189]); 
    assign out[285] = ~(layer_0[7644] ^ layer_0[8363]); 
    assign out[286] = layer_0[9024] & layer_0[6571]; 
    assign out[287] = ~(layer_0[3193] ^ layer_0[10877]); 
    assign out[288] = layer_0[927] ^ layer_0[9735]; 
    assign out[289] = layer_0[10154] ^ layer_0[6653]; 
    assign out[290] = layer_0[1646] ^ layer_0[8573]; 
    assign out[291] = layer_0[8443] ^ layer_0[9945]; 
    assign out[292] = ~(layer_0[10533] & layer_0[7235]); 
    assign out[293] = layer_0[6258] & layer_0[1631]; 
    assign out[294] = layer_0[5497] & layer_0[2760]; 
    assign out[295] = layer_0[5499] & layer_0[3051]; 
    assign out[296] = ~(layer_0[7971] ^ layer_0[9099]); 
    assign out[297] = layer_0[3807] ^ layer_0[1880]; 
    assign out[298] = layer_0[3195] ^ layer_0[4291]; 
    assign out[299] = layer_0[606]; 
    assign out[300] = ~layer_0[2473] | (layer_0[2473] & layer_0[6185]); 
    assign out[301] = ~(layer_0[4382] ^ layer_0[3541]); 
    assign out[302] = ~(layer_0[3499] & layer_0[10396]); 
    assign out[303] = layer_0[6839] ^ layer_0[186]; 
    assign out[304] = layer_0[6649] | layer_0[4882]; 
    assign out[305] = layer_0[6429]; 
    assign out[306] = ~(layer_0[7982] & layer_0[5974]); 
    assign out[307] = layer_0[6401] ^ layer_0[7991]; 
    assign out[308] = layer_0[8895] ^ layer_0[9607]; 
    assign out[309] = layer_0[5285] ^ layer_0[3303]; 
    assign out[310] = layer_0[5156] ^ layer_0[4892]; 
    assign out[311] = ~(layer_0[8701] ^ layer_0[2877]); 
    assign out[312] = ~layer_0[3628] | (layer_0[3628] & layer_0[11904]); 
    assign out[313] = ~(layer_0[5697] ^ layer_0[10591]); 
    assign out[314] = ~(layer_0[9765] ^ layer_0[6]); 
    assign out[315] = ~(layer_0[6227] | layer_0[6436]); 
    assign out[316] = ~(layer_0[9426] & layer_0[976]); 
    assign out[317] = ~(layer_0[4773] ^ layer_0[7881]); 
    assign out[318] = layer_0[8552] ^ layer_0[6226]; 
    assign out[319] = layer_0[2519] & ~layer_0[5989]; 
    assign out[320] = ~(layer_0[8119] ^ layer_0[11634]); 
    assign out[321] = ~layer_0[10602]; 
    assign out[322] = ~(layer_0[7613] & layer_0[4054]); 
    assign out[323] = ~(layer_0[2231] ^ layer_0[6355]); 
    assign out[324] = layer_0[6560]; 
    assign out[325] = layer_0[8480] ^ layer_0[6513]; 
    assign out[326] = ~layer_0[6274]; 
    assign out[327] = layer_0[4718] & ~layer_0[1368]; 
    assign out[328] = layer_0[7490] ^ layer_0[5321]; 
    assign out[329] = ~layer_0[471] | (layer_0[6840] & layer_0[471]); 
    assign out[330] = layer_0[2168] | layer_0[9436]; 
    assign out[331] = ~layer_0[5465] | (layer_0[3472] & layer_0[5465]); 
    assign out[332] = ~(layer_0[6048] ^ layer_0[1429]); 
    assign out[333] = layer_0[2103] ^ layer_0[9074]; 
    assign out[334] = ~(layer_0[11155] ^ layer_0[3330]); 
    assign out[335] = ~layer_0[7520]; 
    assign out[336] = layer_0[1987] ^ layer_0[8296]; 
    assign out[337] = layer_0[10738] ^ layer_0[72]; 
    assign out[338] = layer_0[10321] ^ layer_0[11925]; 
    assign out[339] = ~layer_0[6981]; 
    assign out[340] = ~(layer_0[6071] ^ layer_0[3635]); 
    assign out[341] = ~(layer_0[7107] ^ layer_0[11061]); 
    assign out[342] = ~(layer_0[9736] ^ layer_0[7854]); 
    assign out[343] = ~layer_0[5517] | (layer_0[5517] & layer_0[1025]); 
    assign out[344] = ~(layer_0[9015] ^ layer_0[11071]); 
    assign out[345] = ~(layer_0[11433] ^ layer_0[5348]); 
    assign out[346] = ~layer_0[10215]; 
    assign out[347] = layer_0[868] ^ layer_0[8203]; 
    assign out[348] = layer_0[9397] & layer_0[10697]; 
    assign out[349] = ~(layer_0[11662] ^ layer_0[9838]); 
    assign out[350] = layer_0[8804] ^ layer_0[9575]; 
    assign out[351] = ~(layer_0[2471] ^ layer_0[9259]); 
    assign out[352] = ~(layer_0[4052] ^ layer_0[11098]); 
    assign out[353] = layer_0[7952] & ~layer_0[5002]; 
    assign out[354] = layer_0[3676] ^ layer_0[762]; 
    assign out[355] = ~(layer_0[11184] ^ layer_0[1269]); 
    assign out[356] = layer_0[2532] ^ layer_0[2485]; 
    assign out[357] = ~(layer_0[4995] | layer_0[7972]); 
    assign out[358] = layer_0[3379] ^ layer_0[599]; 
    assign out[359] = ~(layer_0[1730] ^ layer_0[4818]); 
    assign out[360] = layer_0[6590] & layer_0[7148]; 
    assign out[361] = layer_0[295] & layer_0[2548]; 
    assign out[362] = layer_0[9465] ^ layer_0[8656]; 
    assign out[363] = layer_0[5210] & ~layer_0[9616]; 
    assign out[364] = ~layer_0[11325] | (layer_0[9324] & layer_0[11325]); 
    assign out[365] = ~(layer_0[2463] | layer_0[7196]); 
    assign out[366] = ~layer_0[233]; 
    assign out[367] = layer_0[4261] ^ layer_0[673]; 
    assign out[368] = ~(layer_0[3580] ^ layer_0[7]); 
    assign out[369] = ~layer_0[11249]; 
    assign out[370] = ~(layer_0[810] ^ layer_0[6076]); 
    assign out[371] = layer_0[664] ^ layer_0[1314]; 
    assign out[372] = ~(layer_0[4127] & layer_0[9373]); 
    assign out[373] = ~(layer_0[1993] ^ layer_0[5396]); 
    assign out[374] = layer_0[6090] ^ layer_0[4978]; 
    assign out[375] = ~(layer_0[11640] ^ layer_0[8717]); 
    assign out[376] = layer_0[2245]; 
    assign out[377] = layer_0[2781] ^ layer_0[1407]; 
    assign out[378] = layer_0[5780]; 
    assign out[379] = ~layer_0[1037]; 
    assign out[380] = ~(layer_0[10960] ^ layer_0[2252]); 
    assign out[381] = ~(layer_0[7665] | layer_0[11884]); 
    assign out[382] = layer_0[5506] ^ layer_0[6848]; 
    assign out[383] = layer_0[7542] ^ layer_0[4133]; 
    assign out[384] = layer_0[10484] ^ layer_0[8622]; 
    assign out[385] = ~(layer_0[10856] ^ layer_0[944]); 
    assign out[386] = layer_0[990] ^ layer_0[7917]; 
    assign out[387] = ~(layer_0[4153] & layer_0[827]); 
    assign out[388] = layer_0[3966] ^ layer_0[3707]; 
    assign out[389] = layer_0[11967] & ~layer_0[265]; 
    assign out[390] = layer_0[6089]; 
    assign out[391] = layer_0[6902] ^ layer_0[2795]; 
    assign out[392] = layer_0[3979] ^ layer_0[4589]; 
    assign out[393] = ~(layer_0[9647] & layer_0[11952]); 
    assign out[394] = layer_0[6577] ^ layer_0[6749]; 
    assign out[395] = layer_0[11490] ^ layer_0[10838]; 
    assign out[396] = ~(layer_0[7928] ^ layer_0[10077]); 
    assign out[397] = ~layer_0[2113]; 
    assign out[398] = layer_0[8760]; 
    assign out[399] = ~(layer_0[6539] ^ layer_0[1994]); 
    assign out[400] = layer_0[6167] ^ layer_0[10096]; 
    assign out[401] = layer_0[3805] ^ layer_0[6535]; 
    assign out[402] = layer_0[296] ^ layer_0[11652]; 
    assign out[403] = layer_0[9859] ^ layer_0[9445]; 
    assign out[404] = ~(layer_0[9610] ^ layer_0[7747]); 
    assign out[405] = ~(layer_0[1830] & layer_0[7994]); 
    assign out[406] = ~(layer_0[10625] ^ layer_0[2606]); 
    assign out[407] = layer_0[9502] | layer_0[11801]; 
    assign out[408] = layer_0[2328] ^ layer_0[5179]; 
    assign out[409] = layer_0[1487] ^ layer_0[7214]; 
    assign out[410] = layer_0[9164] & layer_0[4696]; 
    assign out[411] = layer_0[34] & ~layer_0[6600]; 
    assign out[412] = layer_0[2089]; 
    assign out[413] = ~(layer_0[3198] ^ layer_0[5608]); 
    assign out[414] = ~layer_0[1057] | (layer_0[8672] & layer_0[1057]); 
    assign out[415] = layer_0[3208] ^ layer_0[785]; 
    assign out[416] = ~layer_0[9824]; 
    assign out[417] = ~layer_0[2250]; 
    assign out[418] = ~(layer_0[9784] ^ layer_0[2264]); 
    assign out[419] = ~(layer_0[1716] ^ layer_0[10264]); 
    assign out[420] = layer_0[5903] ^ layer_0[6218]; 
    assign out[421] = ~(layer_0[690] ^ layer_0[361]); 
    assign out[422] = layer_0[1273] | layer_0[238]; 
    assign out[423] = layer_0[5071]; 
    assign out[424] = layer_0[4142] & ~layer_0[2281]; 
    assign out[425] = layer_0[8110] ^ layer_0[5542]; 
    assign out[426] = ~(layer_0[1417] ^ layer_0[10471]); 
    assign out[427] = layer_0[10461] ^ layer_0[5081]; 
    assign out[428] = layer_0[553] ^ layer_0[223]; 
    assign out[429] = layer_0[10052] ^ layer_0[1235]; 
    assign out[430] = layer_0[8692] & ~layer_0[4648]; 
    assign out[431] = layer_0[10600] & ~layer_0[495]; 
    assign out[432] = layer_0[7464] & layer_0[3797]; 
    assign out[433] = layer_0[2696] ^ layer_0[5174]; 
    assign out[434] = layer_0[11143] ^ layer_0[1590]; 
    assign out[435] = layer_0[2083] ^ layer_0[3271]; 
    assign out[436] = layer_0[10203] ^ layer_0[6669]; 
    assign out[437] = layer_0[2024] & layer_0[336]; 
    assign out[438] = ~(layer_0[10668] & layer_0[1761]); 
    assign out[439] = ~layer_0[4712] | (layer_0[4712] & layer_0[2020]); 
    assign out[440] = layer_0[7057] ^ layer_0[7652]; 
    assign out[441] = ~(layer_0[4296] | layer_0[9469]); 
    assign out[442] = layer_0[4394]; 
    assign out[443] = layer_0[1591] ^ layer_0[5703]; 
    assign out[444] = layer_0[5835] ^ layer_0[11777]; 
    assign out[445] = ~layer_0[5562]; 
    assign out[446] = ~(layer_0[8272] ^ layer_0[297]); 
    assign out[447] = layer_0[7082] ^ layer_0[9084]; 
    assign out[448] = layer_0[8454] ^ layer_0[85]; 
    assign out[449] = ~(layer_0[3132] & layer_0[3571]); 
    assign out[450] = ~layer_0[6680] | (layer_0[1195] & layer_0[6680]); 
    assign out[451] = ~layer_0[8253] | (layer_0[4344] & layer_0[8253]); 
    assign out[452] = ~layer_0[2207]; 
    assign out[453] = ~(layer_0[8144] ^ layer_0[7358]); 
    assign out[454] = ~(layer_0[3562] | layer_0[10225]); 
    assign out[455] = ~(layer_0[2948] ^ layer_0[9097]); 
    assign out[456] = ~layer_0[3233]; 
    assign out[457] = ~(layer_0[5867] ^ layer_0[8965]); 
    assign out[458] = ~layer_0[6761] | (layer_0[4919] & layer_0[6761]); 
    assign out[459] = layer_0[1589]; 
    assign out[460] = layer_0[1173] ^ layer_0[5655]; 
    assign out[461] = ~(layer_0[10233] ^ layer_0[60]); 
    assign out[462] = layer_0[7714]; 
    assign out[463] = layer_0[2220] ^ layer_0[4761]; 
    assign out[464] = layer_0[8469]; 
    assign out[465] = layer_0[10318] & ~layer_0[6209]; 
    assign out[466] = layer_0[11168] ^ layer_0[9328]; 
    assign out[467] = ~layer_0[859]; 
    assign out[468] = ~layer_0[9928] | (layer_0[9928] & layer_0[8936]); 
    assign out[469] = layer_0[9204] ^ layer_0[5031]; 
    assign out[470] = ~(layer_0[5262] | layer_0[1180]); 
    assign out[471] = ~layer_0[2988]; 
    assign out[472] = layer_0[11555] ^ layer_0[5898]; 
    assign out[473] = ~layer_0[10994] | (layer_0[1856] & layer_0[10994]); 
    assign out[474] = layer_0[11388] ^ layer_0[3929]; 
    assign out[475] = layer_0[7173] & ~layer_0[9724]; 
    assign out[476] = layer_0[6490]; 
    assign out[477] = ~(layer_0[6743] ^ layer_0[11701]); 
    assign out[478] = ~(layer_0[299] ^ layer_0[7335]); 
    assign out[479] = layer_0[6511] & layer_0[6148]; 
    assign out[480] = layer_0[4920] ^ layer_0[5483]; 
    assign out[481] = ~layer_0[2164] | (layer_0[2164] & layer_0[10946]); 
    assign out[482] = layer_0[6009]; 
    assign out[483] = layer_0[1838] ^ layer_0[6339]; 
    assign out[484] = ~(layer_0[6500] ^ layer_0[2612]); 
    assign out[485] = layer_0[9629]; 
    assign out[486] = layer_0[2193] & ~layer_0[6631]; 
    assign out[487] = ~layer_0[10911]; 
    assign out[488] = ~(layer_0[6404] & layer_0[10046]); 
    assign out[489] = layer_0[9932] & layer_0[8108]; 
    assign out[490] = ~(layer_0[11400] ^ layer_0[10987]); 
    assign out[491] = ~layer_0[1952] | (layer_0[1952] & layer_0[1438]); 
    assign out[492] = layer_0[9288] ^ layer_0[7482]; 
    assign out[493] = layer_0[6527] ^ layer_0[914]; 
    assign out[494] = ~(layer_0[2993] ^ layer_0[108]); 
    assign out[495] = ~layer_0[1804]; 
    assign out[496] = layer_0[1138] ^ layer_0[8524]; 
    assign out[497] = ~layer_0[11708] | (layer_0[11708] & layer_0[3047]); 
    assign out[498] = ~(layer_0[463] ^ layer_0[1067]); 
    assign out[499] = layer_0[7900] & ~layer_0[936]; 
    assign out[500] = ~(layer_0[11236] ^ layer_0[5161]); 
    assign out[501] = layer_0[3813] & ~layer_0[11908]; 
    assign out[502] = layer_0[6480] | layer_0[9461]; 
    assign out[503] = layer_0[6437] ^ layer_0[4544]; 
    assign out[504] = layer_0[9550] & ~layer_0[11003]; 
    assign out[505] = ~(layer_0[6750] ^ layer_0[6746]); 
    assign out[506] = layer_0[5799]; 
    assign out[507] = layer_0[11142] ^ layer_0[9116]; 
    assign out[508] = layer_0[4243] ^ layer_0[9977]; 
    assign out[509] = ~(layer_0[11429] ^ layer_0[9177]); 
    assign out[510] = ~layer_0[6338] | (layer_0[6338] & layer_0[4207]); 
    assign out[511] = ~(layer_0[5602] & layer_0[185]); 
    assign out[512] = ~layer_0[6274] | (layer_0[6274] & layer_0[10755]); 
    assign out[513] = layer_0[9141] ^ layer_0[2520]; 
    assign out[514] = ~(layer_0[11451] ^ layer_0[348]); 
    assign out[515] = ~layer_0[7455] | (layer_0[8877] & layer_0[7455]); 
    assign out[516] = layer_0[2918] & layer_0[3839]; 
    assign out[517] = ~(layer_0[783] ^ layer_0[6597]); 
    assign out[518] = layer_0[2233] & layer_0[7996]; 
    assign out[519] = layer_0[3376] ^ layer_0[787]; 
    assign out[520] = layer_0[11944] ^ layer_0[6706]; 
    assign out[521] = ~(layer_0[5071] ^ layer_0[642]); 
    assign out[522] = layer_0[1461] ^ layer_0[10665]; 
    assign out[523] = ~layer_0[1430] | (layer_0[1430] & layer_0[8287]); 
    assign out[524] = ~(layer_0[10803] ^ layer_0[3969]); 
    assign out[525] = layer_0[4875] ^ layer_0[1901]; 
    assign out[526] = layer_0[6514] ^ layer_0[771]; 
    assign out[527] = layer_0[7274]; 
    assign out[528] = layer_0[1462] ^ layer_0[9692]; 
    assign out[529] = ~layer_0[1353]; 
    assign out[530] = ~layer_0[3836]; 
    assign out[531] = layer_0[11715] ^ layer_0[922]; 
    assign out[532] = ~(layer_0[6629] ^ layer_0[11897]); 
    assign out[533] = ~(layer_0[1821] & layer_0[10723]); 
    assign out[534] = ~(layer_0[6206] ^ layer_0[8535]); 
    assign out[535] = ~(layer_0[4517] ^ layer_0[10888]); 
    assign out[536] = layer_0[7856] & ~layer_0[8165]; 
    assign out[537] = layer_0[3678] & ~layer_0[3446]; 
    assign out[538] = ~(layer_0[5219] ^ layer_0[10403]); 
    assign out[539] = ~(layer_0[1507] ^ layer_0[11074]); 
    assign out[540] = layer_0[4079] ^ layer_0[6937]; 
    assign out[541] = ~(layer_0[9892] ^ layer_0[5337]); 
    assign out[542] = layer_0[7820] & layer_0[1150]; 
    assign out[543] = layer_0[4263] ^ layer_0[7087]; 
    assign out[544] = layer_0[8229] & ~layer_0[1299]; 
    assign out[545] = ~(layer_0[4860] ^ layer_0[4509]); 
    assign out[546] = ~layer_0[1100] | (layer_0[1100] & layer_0[1280]); 
    assign out[547] = layer_0[4001] ^ layer_0[1897]; 
    assign out[548] = layer_0[7826] ^ layer_0[2126]; 
    assign out[549] = ~(layer_0[8403] ^ layer_0[3801]); 
    assign out[550] = layer_0[191] & layer_0[7492]; 
    assign out[551] = ~layer_0[1378]; 
    assign out[552] = ~(layer_0[9190] ^ layer_0[2574]); 
    assign out[553] = layer_0[6953]; 
    assign out[554] = layer_0[10348] ^ layer_0[6650]; 
    assign out[555] = layer_0[10460] ^ layer_0[2819]; 
    assign out[556] = layer_0[7211] ^ layer_0[299]; 
    assign out[557] = ~layer_0[10947] | (layer_0[10947] & layer_0[136]); 
    assign out[558] = ~(layer_0[3645] ^ layer_0[5211]); 
    assign out[559] = ~(layer_0[8887] ^ layer_0[4865]); 
    assign out[560] = layer_0[1077] | layer_0[2911]; 
    assign out[561] = layer_0[7755] ^ layer_0[11537]; 
    assign out[562] = layer_0[10937] ^ layer_0[9684]; 
    assign out[563] = layer_0[4058] ^ layer_0[7586]; 
    assign out[564] = layer_0[10497] & layer_0[10261]; 
    assign out[565] = layer_0[7792] ^ layer_0[11250]; 
    assign out[566] = layer_0[5777] ^ layer_0[3505]; 
    assign out[567] = layer_0[7794] ^ layer_0[11760]; 
    assign out[568] = layer_0[8640] & layer_0[245]; 
    assign out[569] = layer_0[2570] & layer_0[4788]; 
    assign out[570] = layer_0[2865] ^ layer_0[7642]; 
    assign out[571] = ~(layer_0[11392] ^ layer_0[4144]); 
    assign out[572] = layer_0[686] & layer_0[7926]; 
    assign out[573] = ~layer_0[7901] | (layer_0[8406] & layer_0[7901]); 
    assign out[574] = layer_0[10883] ^ layer_0[6542]; 
    assign out[575] = layer_0[7709] & layer_0[8947]; 
    assign out[576] = layer_0[1001] ^ layer_0[5492]; 
    assign out[577] = layer_0[8482] ^ layer_0[8420]; 
    assign out[578] = layer_0[3743] & ~layer_0[7494]; 
    assign out[579] = ~layer_0[10422]; 
    assign out[580] = layer_0[3959] | layer_0[1443]; 
    assign out[581] = ~(layer_0[9763] ^ layer_0[912]); 
    assign out[582] = layer_0[3524] ^ layer_0[6586]; 
    assign out[583] = layer_0[7451] ^ layer_0[284]; 
    assign out[584] = ~(layer_0[3758] ^ layer_0[3612]); 
    assign out[585] = layer_0[3932] ^ layer_0[8816]; 
    assign out[586] = ~(layer_0[5920] ^ layer_0[2362]); 
    assign out[587] = ~layer_0[9568] | (layer_0[6830] & layer_0[9568]); 
    assign out[588] = layer_0[2088]; 
    assign out[589] = layer_0[6329] ^ layer_0[2331]; 
    assign out[590] = layer_0[1760] ^ layer_0[11078]; 
    assign out[591] = layer_0[5473] ^ layer_0[8718]; 
    assign out[592] = layer_0[8601]; 
    assign out[593] = ~(layer_0[2817] ^ layer_0[522]); 
    assign out[594] = ~(layer_0[11953] ^ layer_0[1445]); 
    assign out[595] = ~layer_0[4395] | (layer_0[4395] & layer_0[8362]); 
    assign out[596] = layer_0[729] ^ layer_0[7958]; 
    assign out[597] = layer_0[7252] & ~layer_0[2432]; 
    assign out[598] = layer_0[4577]; 
    assign out[599] = layer_0[4800] ^ layer_0[2121]; 
    assign out[600] = ~(layer_0[1938] ^ layer_0[9550]); 
    assign out[601] = ~(layer_0[5830] & layer_0[10571]); 
    assign out[602] = layer_0[7997] ^ layer_0[5165]; 
    assign out[603] = ~(layer_0[10407] ^ layer_0[1267]); 
    assign out[604] = layer_0[9565]; 
    assign out[605] = ~layer_0[575] | (layer_0[575] & layer_0[1674]); 
    assign out[606] = ~layer_0[10759]; 
    assign out[607] = ~(layer_0[5443] ^ layer_0[11216]); 
    assign out[608] = layer_0[5610] ^ layer_0[2363]; 
    assign out[609] = ~(layer_0[6990] ^ layer_0[10481]); 
    assign out[610] = layer_0[4393] & layer_0[2968]; 
    assign out[611] = layer_0[8375] ^ layer_0[10375]; 
    assign out[612] = ~(layer_0[11824] ^ layer_0[10223]); 
    assign out[613] = ~(layer_0[5433] ^ layer_0[7573]); 
    assign out[614] = layer_0[10075] ^ layer_0[11967]; 
    assign out[615] = layer_0[1499]; 
    assign out[616] = layer_0[836] & ~layer_0[11005]; 
    assign out[617] = layer_0[8965] ^ layer_0[1627]; 
    assign out[618] = layer_0[412] ^ layer_0[9396]; 
    assign out[619] = ~layer_0[5688] | (layer_0[9532] & layer_0[5688]); 
    assign out[620] = layer_0[10901]; 
    assign out[621] = layer_0[9519] ^ layer_0[1922]; 
    assign out[622] = ~(layer_0[1871] & layer_0[8603]); 
    assign out[623] = ~(layer_0[970] ^ layer_0[9752]); 
    assign out[624] = ~(layer_0[11593] ^ layer_0[5139]); 
    assign out[625] = ~(layer_0[8198] | layer_0[11877]); 
    assign out[626] = layer_0[11890] & layer_0[11554]; 
    assign out[627] = ~(layer_0[10350] ^ layer_0[6985]); 
    assign out[628] = layer_0[8210]; 
    assign out[629] = ~(layer_0[11233] ^ layer_0[10273]); 
    assign out[630] = ~(layer_0[11711] ^ layer_0[3506]); 
    assign out[631] = layer_0[2112] & layer_0[10381]; 
    assign out[632] = layer_0[7949]; 
    assign out[633] = ~layer_0[8677] | (layer_0[8677] & layer_0[7288]); 
    assign out[634] = ~(layer_0[8565] | layer_0[2091]); 
    assign out[635] = layer_0[9759] ^ layer_0[4224]; 
    assign out[636] = ~(layer_0[10208] ^ layer_0[5674]); 
    assign out[637] = ~(layer_0[6950] ^ layer_0[1723]); 
    assign out[638] = ~layer_0[2334] | (layer_0[11935] & layer_0[2334]); 
    assign out[639] = layer_0[9946] & layer_0[3525]; 
    assign out[640] = layer_0[5142] ^ layer_0[8278]; 
    assign out[641] = layer_0[10191]; 
    assign out[642] = ~layer_0[4351] | (layer_0[4351] & layer_0[1214]); 
    assign out[643] = layer_0[2926] & ~layer_0[10412]; 
    assign out[644] = layer_0[8331] ^ layer_0[5567]; 
    assign out[645] = ~(layer_0[8696] ^ layer_0[5319]); 
    assign out[646] = ~(layer_0[5615] ^ layer_0[9823]); 
    assign out[647] = layer_0[9455]; 
    assign out[648] = ~layer_0[11389] | (layer_0[8186] & layer_0[11389]); 
    assign out[649] = ~(layer_0[4972] ^ layer_0[10240]); 
    assign out[650] = layer_0[7460] ^ layer_0[8188]; 
    assign out[651] = layer_0[613] ^ layer_0[8349]; 
    assign out[652] = ~(layer_0[356] ^ layer_0[1568]); 
    assign out[653] = ~layer_0[302]; 
    assign out[654] = layer_0[8020] ^ layer_0[5847]; 
    assign out[655] = layer_0[9588] ^ layer_0[7404]; 
    assign out[656] = layer_0[2358] ^ layer_0[1492]; 
    assign out[657] = layer_0[7304] ^ layer_0[3815]; 
    assign out[658] = ~(layer_0[6948] ^ layer_0[7993]); 
    assign out[659] = layer_0[7364] | layer_0[11416]; 
    assign out[660] = layer_0[3305] ^ layer_0[11870]; 
    assign out[661] = ~layer_0[11626] | (layer_0[11626] & layer_0[7903]); 
    assign out[662] = ~(layer_0[5166] ^ layer_0[393]); 
    assign out[663] = layer_0[11699] ^ layer_0[2955]; 
    assign out[664] = layer_0[3709] ^ layer_0[11354]; 
    assign out[665] = layer_0[7967] & ~layer_0[3136]; 
    assign out[666] = layer_0[5593] & ~layer_0[8098]; 
    assign out[667] = ~(layer_0[8154] ^ layer_0[3690]); 
    assign out[668] = ~(layer_0[888] ^ layer_0[11247]); 
    assign out[669] = layer_0[11466] & ~layer_0[6827]; 
    assign out[670] = ~layer_0[2976]; 
    assign out[671] = layer_0[1506] ^ layer_0[8707]; 
    assign out[672] = ~(layer_0[6862] ^ layer_0[4970]); 
    assign out[673] = ~(layer_0[10731] ^ layer_0[3254]); 
    assign out[674] = layer_0[5664] ^ layer_0[11675]; 
    assign out[675] = layer_0[5196] & ~layer_0[1688]; 
    assign out[676] = layer_0[6458]; 
    assign out[677] = layer_0[604] ^ layer_0[6459]; 
    assign out[678] = ~(layer_0[3045] ^ layer_0[6288]); 
    assign out[679] = layer_0[1567] ^ layer_0[11407]; 
    assign out[680] = layer_0[2972] & ~layer_0[1865]; 
    assign out[681] = layer_0[10260] ^ layer_0[6978]; 
    assign out[682] = ~(layer_0[5527] ^ layer_0[7333]); 
    assign out[683] = layer_0[8209] ^ layer_0[6644]; 
    assign out[684] = layer_0[7074] & ~layer_0[11415]; 
    assign out[685] = layer_0[2242] & ~layer_0[956]; 
    assign out[686] = ~(layer_0[563] ^ layer_0[5163]); 
    assign out[687] = ~(layer_0[7349] ^ layer_0[436]); 
    assign out[688] = layer_0[5324] & ~layer_0[7013]; 
    assign out[689] = ~(layer_0[6219] ^ layer_0[11912]); 
    assign out[690] = ~layer_0[1172] | (layer_0[1172] & layer_0[5537]); 
    assign out[691] = layer_0[8175] ^ layer_0[857]; 
    assign out[692] = ~(layer_0[1206] & layer_0[2831]); 
    assign out[693] = layer_0[83]; 
    assign out[694] = layer_0[10763] & layer_0[10790]; 
    assign out[695] = layer_0[4329] ^ layer_0[8661]; 
    assign out[696] = layer_0[11510] & ~layer_0[659]; 
    assign out[697] = layer_0[665] ^ layer_0[704]; 
    assign out[698] = ~layer_0[3772]; 
    assign out[699] = layer_0[11954] ^ layer_0[2247]; 
    assign out[700] = layer_0[1707] ^ layer_0[2107]; 
    assign out[701] = layer_0[355] & ~layer_0[5489]; 
    assign out[702] = ~layer_0[2263] | (layer_0[8483] & layer_0[2263]); 
    assign out[703] = layer_0[5590]; 
    assign out[704] = ~(layer_0[3273] ^ layer_0[4489]); 
    assign out[705] = layer_0[3486] ^ layer_0[11029]; 
    assign out[706] = ~(layer_0[9014] ^ layer_0[11167]); 
    assign out[707] = layer_0[6174] ^ layer_0[4216]; 
    assign out[708] = ~layer_0[4104] | (layer_0[4104] & layer_0[1109]); 
    assign out[709] = ~(layer_0[10983] ^ layer_0[7602]); 
    assign out[710] = ~(layer_0[9962] & layer_0[5084]); 
    assign out[711] = layer_0[4836] ^ layer_0[7578]; 
    assign out[712] = ~(layer_0[8465] ^ layer_0[8023]); 
    assign out[713] = ~(layer_0[1603] ^ layer_0[4571]); 
    assign out[714] = ~(layer_0[8727] ^ layer_0[9534]); 
    assign out[715] = layer_0[272] ^ layer_0[1124]; 
    assign out[716] = ~(layer_0[7623] ^ layer_0[5401]); 
    assign out[717] = layer_0[5998] ^ layer_0[2321]; 
    assign out[718] = layer_0[10148] ^ layer_0[1518]; 
    assign out[719] = layer_0[5557] & ~layer_0[6442]; 
    assign out[720] = ~(layer_0[1598] ^ layer_0[11609]); 
    assign out[721] = ~(layer_0[2368] | layer_0[1888]); 
    assign out[722] = ~(layer_0[10131] ^ layer_0[780]); 
    assign out[723] = layer_0[8941]; 
    assign out[724] = layer_0[6956]; 
    assign out[725] = layer_0[6178] | layer_0[8724]; 
    assign out[726] = ~layer_0[11207]; 
    assign out[727] = layer_0[7150]; 
    assign out[728] = ~(layer_0[2243] ^ layer_0[9967]); 
    assign out[729] = ~(layer_0[7466] ^ layer_0[6204]); 
    assign out[730] = ~(layer_0[6276] ^ layer_0[6280]); 
    assign out[731] = ~(layer_0[4554] | layer_0[20]); 
    assign out[732] = ~layer_0[446] | (layer_0[1159] & layer_0[446]); 
    assign out[733] = layer_0[9397]; 
    assign out[734] = layer_0[7562]; 
    assign out[735] = layer_0[4340] ^ layer_0[8649]; 
    assign out[736] = layer_0[8180] ^ layer_0[5271]; 
    assign out[737] = ~layer_0[5664]; 
    assign out[738] = layer_0[11023] | layer_0[6172]; 
    assign out[739] = ~(layer_0[1522] ^ layer_0[3738]); 
    assign out[740] = layer_0[2767] ^ layer_0[86]; 
    assign out[741] = layer_0[3978] ^ layer_0[11587]; 
    assign out[742] = layer_0[6118] ^ layer_0[1784]; 
    assign out[743] = ~(layer_0[5241] ^ layer_0[10437]); 
    assign out[744] = layer_0[5685] ^ layer_0[10623]; 
    assign out[745] = layer_0[11177] & ~layer_0[10238]; 
    assign out[746] = ~layer_0[5961] | (layer_0[8584] & layer_0[5961]); 
    assign out[747] = ~(layer_0[4615] | layer_0[6757]); 
    assign out[748] = layer_0[9897] ^ layer_0[7809]; 
    assign out[749] = ~(layer_0[10174] | layer_0[1226]); 
    assign out[750] = ~(layer_0[11678] | layer_0[9487]); 
    assign out[751] = layer_0[5969] ^ layer_0[7708]; 
    assign out[752] = layer_0[127]; 
    assign out[753] = layer_0[1432] & ~layer_0[774]; 
    assign out[754] = ~(layer_0[2751] & layer_0[1184]); 
    assign out[755] = layer_0[11370]; 
    assign out[756] = ~layer_0[8914] | (layer_0[8914] & layer_0[2355]); 
    assign out[757] = ~(layer_0[11759] | layer_0[5012]); 
    assign out[758] = layer_0[6198] ^ layer_0[2795]; 
    assign out[759] = ~(layer_0[11148] & layer_0[2461]); 
    assign out[760] = layer_0[909] & ~layer_0[11654]; 
    assign out[761] = layer_0[8653] ^ layer_0[5256]; 
    assign out[762] = ~(layer_0[4768] ^ layer_0[11321]); 
    assign out[763] = ~(layer_0[3592] | layer_0[1762]); 
    assign out[764] = layer_0[11031]; 
    assign out[765] = ~(layer_0[11067] & layer_0[2697]); 
    assign out[766] = layer_0[6561] ^ layer_0[1717]; 
    assign out[767] = layer_0[6221] & layer_0[466]; 
    assign out[768] = layer_0[7063] & layer_0[8220]; 
    assign out[769] = layer_0[2882] | layer_0[3445]; 
    assign out[770] = ~(layer_0[7056] ^ layer_0[11621]); 
    assign out[771] = layer_0[10965] ^ layer_0[4049]; 
    assign out[772] = ~(layer_0[5728] ^ layer_0[5180]); 
    assign out[773] = ~layer_0[10784]; 
    assign out[774] = layer_0[11487]; 
    assign out[775] = layer_0[4683] ^ layer_0[5840]; 
    assign out[776] = layer_0[3397] & ~layer_0[6283]; 
    assign out[777] = ~(layer_0[9493] ^ layer_0[8443]); 
    assign out[778] = layer_0[760] ^ layer_0[5849]; 
    assign out[779] = layer_0[11789] ^ layer_0[10513]; 
    assign out[780] = layer_0[9899] & ~layer_0[68]; 
    assign out[781] = ~(layer_0[8773] ^ layer_0[10967]); 
    assign out[782] = layer_0[1798] & ~layer_0[11535]; 
    assign out[783] = ~(layer_0[4092] | layer_0[2353]); 
    assign out[784] = layer_0[1632] & ~layer_0[6635]; 
    assign out[785] = ~layer_0[8114] | (layer_0[8114] & layer_0[723]); 
    assign out[786] = layer_0[5662] & layer_0[10526]; 
    assign out[787] = ~layer_0[4008]; 
    assign out[788] = layer_0[3162] & ~layer_0[8620]; 
    assign out[789] = layer_0[8786] ^ layer_0[2543]; 
    assign out[790] = ~(layer_0[10057] & layer_0[6701]); 
    assign out[791] = ~(layer_0[2829] ^ layer_0[5208]); 
    assign out[792] = layer_0[8388] & ~layer_0[70]; 
    assign out[793] = layer_0[1903] ^ layer_0[3590]; 
    assign out[794] = layer_0[7371] ^ layer_0[6931]; 
    assign out[795] = ~(layer_0[10613] ^ layer_0[5888]); 
    assign out[796] = ~layer_0[2094] | (layer_0[3471] & layer_0[2094]); 
    assign out[797] = ~(layer_0[3506] ^ layer_0[2870]); 
    assign out[798] = layer_0[2047] | layer_0[8521]; 
    assign out[799] = layer_0[6369] ^ layer_0[6754]; 
    assign out[800] = layer_0[8562] & ~layer_0[375]; 
    assign out[801] = ~(layer_0[5702] ^ layer_0[1513]); 
    assign out[802] = layer_0[1424] ^ layer_0[4124]; 
    assign out[803] = layer_0[2752] & layer_0[7386]; 
    assign out[804] = ~(layer_0[5277] ^ layer_0[3069]); 
    assign out[805] = ~layer_0[2538]; 
    assign out[806] = ~layer_0[8462] | (layer_0[9929] & layer_0[8462]); 
    assign out[807] = ~(layer_0[6607] ^ layer_0[10716]); 
    assign out[808] = layer_0[10378]; 
    assign out[809] = layer_0[3501] ^ layer_0[1516]; 
    assign out[810] = ~(layer_0[11719] & layer_0[10644]); 
    assign out[811] = ~(layer_0[146] | layer_0[10305]); 
    assign out[812] = layer_0[4198] ^ layer_0[7487]; 
    assign out[813] = layer_0[6488] ^ layer_0[7688]; 
    assign out[814] = ~(layer_0[10007] ^ layer_0[2858]); 
    assign out[815] = layer_0[7424]; 
    assign out[816] = ~(layer_0[9921] | layer_0[2822]); 
    assign out[817] = ~(layer_0[8559] ^ layer_0[8706]); 
    assign out[818] = layer_0[8046] ^ layer_0[4799]; 
    assign out[819] = ~(layer_0[9574] ^ layer_0[2051]); 
    assign out[820] = layer_0[1787] & layer_0[5521]; 
    assign out[821] = ~(layer_0[6877] ^ layer_0[10822]); 
    assign out[822] = layer_0[6894] ^ layer_0[8959]; 
    assign out[823] = layer_0[6849]; 
    assign out[824] = ~(layer_0[9219] | layer_0[5024]); 
    assign out[825] = ~(layer_0[5250] ^ layer_0[1020]); 
    assign out[826] = ~layer_0[3965]; 
    assign out[827] = layer_0[187] & ~layer_0[10083]; 
    assign out[828] = ~layer_0[4813]; 
    assign out[829] = layer_0[9256]; 
    assign out[830] = layer_0[3644] & layer_0[2032]; 
    assign out[831] = ~(layer_0[2990] & layer_0[9773]); 
    assign out[832] = ~(layer_0[5619] ^ layer_0[2675]); 
    assign out[833] = ~layer_0[1065] | (layer_0[1065] & layer_0[4957]); 
    assign out[834] = layer_0[887]; 
    assign out[835] = layer_0[11394]; 
    assign out[836] = layer_0[219] ^ layer_0[6637]; 
    assign out[837] = layer_0[1387] & layer_0[11320]; 
    assign out[838] = ~(layer_0[813] ^ layer_0[2417]); 
    assign out[839] = layer_0[11706] & ~layer_0[595]; 
    assign out[840] = layer_0[4028]; 
    assign out[841] = ~layer_0[5049] | (layer_0[8570] & layer_0[5049]); 
    assign out[842] = layer_0[11558] ^ layer_0[2787]; 
    assign out[843] = layer_0[11228] ^ layer_0[9537]; 
    assign out[844] = layer_0[5909] ^ layer_0[6601]; 
    assign out[845] = layer_0[3630] ^ layer_0[6312]; 
    assign out[846] = layer_0[1541] & ~layer_0[8838]; 
    assign out[847] = ~(layer_0[11691] | layer_0[3117]); 
    assign out[848] = layer_0[10042] ^ layer_0[1819]; 
    assign out[849] = layer_0[3649] & layer_0[7853]; 
    assign out[850] = layer_0[1557] ^ layer_0[10778]; 
    assign out[851] = ~layer_0[10309] | (layer_0[6949] & layer_0[10309]); 
    assign out[852] = ~layer_0[9596] | (layer_0[9596] & layer_0[654]); 
    assign out[853] = ~layer_0[2486]; 
    assign out[854] = layer_0[11677] ^ layer_0[1607]; 
    assign out[855] = layer_0[5915]; 
    assign out[856] = layer_0[578] ^ layer_0[4020]; 
    assign out[857] = layer_0[4193] & ~layer_0[7159]; 
    assign out[858] = ~(layer_0[3768] ^ layer_0[8935]); 
    assign out[859] = layer_0[1996]; 
    assign out[860] = ~(layer_0[4247] ^ layer_0[7635]); 
    assign out[861] = ~layer_0[7203]; 
    assign out[862] = layer_0[1192]; 
    assign out[863] = layer_0[10526]; 
    assign out[864] = ~(layer_0[3399] ^ layer_0[3314]); 
    assign out[865] = layer_0[7265]; 
    assign out[866] = ~layer_0[8407] | (layer_0[4905] & layer_0[8407]); 
    assign out[867] = layer_0[6385]; 
    assign out[868] = ~(layer_0[9544] ^ layer_0[9689]); 
    assign out[869] = ~(layer_0[9470] ^ layer_0[5270]); 
    assign out[870] = layer_0[10549] ^ layer_0[1359]; 
    assign out[871] = ~(layer_0[2283] ^ layer_0[10207]); 
    assign out[872] = ~layer_0[7204]; 
    assign out[873] = layer_0[3039] ^ layer_0[7841]; 
    assign out[874] = layer_0[7652]; 
    assign out[875] = ~layer_0[10819]; 
    assign out[876] = ~layer_0[4780] | (layer_0[4780] & layer_0[9728]); 
    assign out[877] = ~layer_0[4635]; 
    assign out[878] = ~layer_0[4766]; 
    assign out[879] = layer_0[2408] ^ layer_0[11284]; 
    assign out[880] = ~(layer_0[11316] ^ layer_0[3945]); 
    assign out[881] = ~layer_0[3056]; 
    assign out[882] = layer_0[6015] ^ layer_0[2961]; 
    assign out[883] = ~layer_0[5110] | (layer_0[5110] & layer_0[8451]); 
    assign out[884] = layer_0[11208] ^ layer_0[11832]; 
    assign out[885] = layer_0[7137] ^ layer_0[5640]; 
    assign out[886] = layer_0[3849] & layer_0[9514]; 
    assign out[887] = ~layer_0[2528] | (layer_0[9799] & layer_0[2528]); 
    assign out[888] = layer_0[3067] & ~layer_0[8103]; 
    assign out[889] = ~(layer_0[1055] ^ layer_0[6823]); 
    assign out[890] = layer_0[8091]; 
    assign out[891] = layer_0[8221] & ~layer_0[9199]; 
    assign out[892] = layer_0[7827] & layer_0[10962]; 
    assign out[893] = layer_0[5770]; 
    assign out[894] = ~(layer_0[7640] ^ layer_0[7575]); 
    assign out[895] = layer_0[5596]; 
    assign out[896] = ~(layer_0[4277] ^ layer_0[3519]); 
    assign out[897] = layer_0[7718] & ~layer_0[7528]; 
    assign out[898] = layer_0[4456] & layer_0[7828]; 
    assign out[899] = ~layer_0[3166]; 
    assign out[900] = ~(layer_0[10425] ^ layer_0[4232]); 
    assign out[901] = ~(layer_0[2224] ^ layer_0[5753]); 
    assign out[902] = layer_0[10345]; 
    assign out[903] = ~(layer_0[4288] ^ layer_0[10209]); 
    assign out[904] = layer_0[11513] ^ layer_0[8057]; 
    assign out[905] = layer_0[10930] & ~layer_0[2658]; 
    assign out[906] = layer_0[3012]; 
    assign out[907] = layer_0[11656]; 
    assign out[908] = layer_0[8398]; 
    assign out[909] = layer_0[6470] ^ layer_0[1858]; 
    assign out[910] = ~(layer_0[2589] ^ layer_0[3943]); 
    assign out[911] = ~(layer_0[2158] & layer_0[4526]); 
    assign out[912] = layer_0[3515] ^ layer_0[2576]; 
    assign out[913] = ~layer_0[1695] | (layer_0[31] & layer_0[1695]); 
    assign out[914] = layer_0[5260] & layer_0[7319]; 
    assign out[915] = layer_0[2178] & ~layer_0[10234]; 
    assign out[916] = layer_0[5657]; 
    assign out[917] = layer_0[4179] ^ layer_0[9914]; 
    assign out[918] = layer_0[5733]; 
    assign out[919] = layer_0[3100] & ~layer_0[3213]; 
    assign out[920] = layer_0[5875] | layer_0[2483]; 
    assign out[921] = layer_0[11015]; 
    assign out[922] = layer_0[963]; 
    assign out[923] = ~(layer_0[7438] & layer_0[8246]); 
    assign out[924] = layer_0[3859]; 
    assign out[925] = ~layer_0[3742]; 
    assign out[926] = layer_0[5612] ^ layer_0[5797]; 
    assign out[927] = ~(layer_0[796] ^ layer_0[343]); 
    assign out[928] = layer_0[1309] & layer_0[1909]; 
    assign out[929] = ~(layer_0[992] & layer_0[11127]); 
    assign out[930] = layer_0[9474]; 
    assign out[931] = ~layer_0[4812]; 
    assign out[932] = ~(layer_0[5579] ^ layer_0[8138]); 
    assign out[933] = ~(layer_0[1644] ^ layer_0[11384]); 
    assign out[934] = ~(layer_0[11768] | layer_0[9778]); 
    assign out[935] = ~(layer_0[10206] ^ layer_0[88]); 
    assign out[936] = layer_0[2577]; 
    assign out[937] = layer_0[7108] ^ layer_0[9481]; 
    assign out[938] = layer_0[10387] ^ layer_0[2810]; 
    assign out[939] = layer_0[3191] ^ layer_0[3685]; 
    assign out[940] = layer_0[2027] & layer_0[2991]; 
    assign out[941] = layer_0[9241] ^ layer_0[8606]; 
    assign out[942] = layer_0[5871] | layer_0[6482]; 
    assign out[943] = layer_0[2588] & ~layer_0[7210]; 
    assign out[944] = layer_0[8986] ^ layer_0[4697]; 
    assign out[945] = layer_0[1419]; 
    assign out[946] = layer_0[320] & ~layer_0[5784]; 
    assign out[947] = ~layer_0[1972]; 
    assign out[948] = ~(layer_0[10899] ^ layer_0[4191]); 
    assign out[949] = layer_0[439] ^ layer_0[7436]; 
    assign out[950] = layer_0[329] ^ layer_0[8078]; 
    assign out[951] = layer_0[10157] ^ layer_0[9561]; 
    assign out[952] = layer_0[43]; 
    assign out[953] = layer_0[10596] & ~layer_0[4732]; 
    assign out[954] = layer_0[9421] & ~layer_0[11712]; 
    assign out[955] = ~(layer_0[6593] ^ layer_0[7034]); 
    assign out[956] = layer_0[9302] & ~layer_0[1379]; 
    assign out[957] = layer_0[10704] ^ layer_0[4218]; 
    assign out[958] = layer_0[1241] & ~layer_0[764]; 
    assign out[959] = ~layer_0[4634] | (layer_0[4634] & layer_0[7041]); 
    assign out[960] = ~(layer_0[1697] ^ layer_0[853]); 
    assign out[961] = layer_0[10133] ^ layer_0[500]; 
    assign out[962] = ~(layer_0[7842] ^ layer_0[10048]); 
    assign out[963] = layer_0[9683] | layer_0[4838]; 
    assign out[964] = layer_0[3055] & ~layer_0[7622]; 
    assign out[965] = layer_0[6353] ^ layer_0[6424]; 
    assign out[966] = ~(layer_0[1061] ^ layer_0[10464]); 
    assign out[967] = ~(layer_0[10651] ^ layer_0[8281]); 
    assign out[968] = ~layer_0[2814]; 
    assign out[969] = ~(layer_0[3317] ^ layer_0[8429]); 
    assign out[970] = layer_0[6635]; 
    assign out[971] = layer_0[7886] ^ layer_0[910]; 
    assign out[972] = ~(layer_0[8874] ^ layer_0[3485]); 
    assign out[973] = ~layer_0[11821] | (layer_0[11821] & layer_0[7851]); 
    assign out[974] = layer_0[10241] & layer_0[10040]; 
    assign out[975] = layer_0[2313]; 
    assign out[976] = layer_0[9448] & layer_0[8906]; 
    assign out[977] = layer_0[6107] & ~layer_0[1785]; 
    assign out[978] = layer_0[4442] ^ layer_0[1444]; 
    assign out[979] = layer_0[11902]; 
    assign out[980] = ~(layer_0[11800] ^ layer_0[6738]); 
    assign out[981] = layer_0[4125] ^ layer_0[2058]; 
    assign out[982] = ~(layer_0[794] ^ layer_0[527]); 
    assign out[983] = ~layer_0[7700]; 
    assign out[984] = layer_0[10509] & ~layer_0[4158]; 
    assign out[985] = ~(layer_0[3732] ^ layer_0[11501]); 
    assign out[986] = ~(layer_0[5642] ^ layer_0[266]); 
    assign out[987] = ~(layer_0[7847] ^ layer_0[5099]); 
    assign out[988] = layer_0[6559] & ~layer_0[9668]; 
    assign out[989] = ~layer_0[2526]; 
    assign out[990] = ~layer_0[7952]; 
    assign out[991] = layer_0[4332] ^ layer_0[2871]; 
    assign out[992] = layer_0[3713] ^ layer_0[10554]; 
    assign out[993] = layer_0[6780] & ~layer_0[2554]; 
    assign out[994] = ~(layer_0[10900] ^ layer_0[6718]); 
    assign out[995] = layer_0[3911] & ~layer_0[445]; 
    assign out[996] = layer_0[11784] ^ layer_0[5157]; 
    assign out[997] = layer_0[5692] & layer_0[10152]; 
    assign out[998] = ~layer_0[9887]; 
    assign out[999] = ~layer_0[3971] | (layer_0[3971] & layer_0[4767]); 
    assign out[1000] = layer_0[7517] ^ layer_0[3143]; 
    assign out[1001] = ~layer_0[8385]; 
    assign out[1002] = layer_0[3345] & layer_0[4825]; 
    assign out[1003] = layer_0[9339] ^ layer_0[9087]; 
    assign out[1004] = ~layer_0[2613] | (layer_0[6181] & layer_0[2613]); 
    assign out[1005] = ~(layer_0[7858] ^ layer_0[3972]); 
    assign out[1006] = ~layer_0[1264]; 
    assign out[1007] = layer_0[4802]; 
    assign out[1008] = layer_0[10006] | layer_0[197]; 
    assign out[1009] = layer_0[2559]; 
    assign out[1010] = layer_0[6807] ^ layer_0[4511]; 
    assign out[1011] = ~(layer_0[9609] ^ layer_0[468]); 
    assign out[1012] = ~(layer_0[6352] | layer_0[5763]); 
    assign out[1013] = layer_0[2004] ^ layer_0[3051]; 
    assign out[1014] = ~layer_0[8564]; 
    assign out[1015] = layer_0[1449]; 
    assign out[1016] = ~(layer_0[8153] ^ layer_0[8987]); 
    assign out[1017] = ~layer_0[6035] | (layer_0[6035] & layer_0[9663]); 
    assign out[1018] = layer_0[6080] ^ layer_0[1365]; 
    assign out[1019] = ~layer_0[10227] | (layer_0[4233] & layer_0[10227]); 
    assign out[1020] = ~(layer_0[473] & layer_0[7023]); 
    assign out[1021] = layer_0[4584]; 
    assign out[1022] = layer_0[8170] & ~layer_0[9539]; 
    assign out[1023] = ~layer_0[228]; 
    assign out[1024] = ~layer_0[10710]; 
    assign out[1025] = layer_0[7307] ^ layer_0[1561]; 
    assign out[1026] = layer_0[667] ^ layer_0[6397]; 
    assign out[1027] = ~layer_0[10192]; 
    assign out[1028] = layer_0[7405] & ~layer_0[8075]; 
    assign out[1029] = layer_0[6019] & layer_0[7158]; 
    assign out[1030] = ~layer_0[3500]; 
    assign out[1031] = layer_0[2611] ^ layer_0[6307]; 
    assign out[1032] = layer_0[11222] & ~layer_0[9239]; 
    assign out[1033] = layer_0[2322] ^ layer_0[11176]; 
    assign out[1034] = ~(layer_0[11050] ^ layer_0[587]); 
    assign out[1035] = ~(layer_0[11334] ^ layer_0[3141]); 
    assign out[1036] = layer_0[2994]; 
    assign out[1037] = layer_0[4101] & ~layer_0[6526]; 
    assign out[1038] = layer_0[8380]; 
    assign out[1039] = layer_0[10972] & ~layer_0[2301]; 
    assign out[1040] = layer_0[6774] ^ layer_0[5932]; 
    assign out[1041] = layer_0[11685] & layer_0[10833]; 
    assign out[1042] = layer_0[2680] ^ layer_0[657]; 
    assign out[1043] = ~(layer_0[7280] ^ layer_0[5620]); 
    assign out[1044] = layer_0[2779] & layer_0[1135]; 
    assign out[1045] = layer_0[10959] ^ layer_0[10201]; 
    assign out[1046] = layer_0[5441] ^ layer_0[11595]; 
    assign out[1047] = ~(layer_0[2710] & layer_0[9093]); 
    assign out[1048] = ~(layer_0[8183] ^ layer_0[7566]); 
    assign out[1049] = layer_0[8422] | layer_0[358]; 
    assign out[1050] = ~(layer_0[11872] | layer_0[1297]); 
    assign out[1051] = ~(layer_0[5248] ^ layer_0[3300]); 
    assign out[1052] = layer_0[2637] & ~layer_0[10315]; 
    assign out[1053] = layer_0[11614] & layer_0[9709]; 
    assign out[1054] = layer_0[1535]; 
    assign out[1055] = ~layer_0[2148]; 
    assign out[1056] = ~(layer_0[9998] ^ layer_0[7989]); 
    assign out[1057] = ~layer_0[6703]; 
    assign out[1058] = layer_0[4762] & layer_0[3590]; 
    assign out[1059] = ~(layer_0[2284] ^ layer_0[2808]); 
    assign out[1060] = ~(layer_0[7564] ^ layer_0[3013]); 
    assign out[1061] = layer_0[1732] & ~layer_0[2901]; 
    assign out[1062] = ~layer_0[10028]; 
    assign out[1063] = ~layer_0[10936]; 
    assign out[1064] = ~(layer_0[7045] ^ layer_0[9299]); 
    assign out[1065] = ~(layer_0[9476] ^ layer_0[972]); 
    assign out[1066] = ~(layer_0[8214] ^ layer_0[6917]); 
    assign out[1067] = layer_0[3335] ^ layer_0[11817]; 
    assign out[1068] = ~layer_0[8342]; 
    assign out[1069] = layer_0[10183]; 
    assign out[1070] = ~(layer_0[11057] ^ layer_0[10292]); 
    assign out[1071] = layer_0[2096] ^ layer_0[9162]; 
    assign out[1072] = ~(layer_0[7290] ^ layer_0[1348]); 
    assign out[1073] = layer_0[10205] ^ layer_0[9285]; 
    assign out[1074] = ~(layer_0[3142] | layer_0[7126]); 
    assign out[1075] = layer_0[9852] & layer_0[6402]; 
    assign out[1076] = ~(layer_0[2109] | layer_0[2403]); 
    assign out[1077] = ~(layer_0[1179] ^ layer_0[4267]); 
    assign out[1078] = ~(layer_0[2828] ^ layer_0[6220]); 
    assign out[1079] = layer_0[8506] & layer_0[1307]; 
    assign out[1080] = layer_0[6495] ^ layer_0[8606]; 
    assign out[1081] = ~(layer_0[10715] ^ layer_0[11903]); 
    assign out[1082] = layer_0[685]; 
    assign out[1083] = layer_0[4627] & ~layer_0[11840]; 
    assign out[1084] = layer_0[1932] & layer_0[3843]; 
    assign out[1085] = layer_0[10726] & ~layer_0[1284]; 
    assign out[1086] = ~layer_0[8445]; 
    assign out[1087] = layer_0[7412] ^ layer_0[7479]; 
    assign out[1088] = ~(layer_0[11358] ^ layer_0[5376]); 
    assign out[1089] = layer_0[8267] ^ layer_0[7712]; 
    assign out[1090] = layer_0[11702] ^ layer_0[1795]; 
    assign out[1091] = ~layer_0[1108] | (layer_0[371] & layer_0[1108]); 
    assign out[1092] = layer_0[9183] & layer_0[5094]; 
    assign out[1093] = ~(layer_0[2410] ^ layer_0[10816]); 
    assign out[1094] = ~(layer_0[5942] | layer_0[10376]); 
    assign out[1095] = layer_0[2196] ^ layer_0[9195]; 
    assign out[1096] = layer_0[1374] ^ layer_0[5289]; 
    assign out[1097] = layer_0[367] ^ layer_0[11990]; 
    assign out[1098] = ~layer_0[7462] | (layer_0[5604] & layer_0[7462]); 
    assign out[1099] = layer_0[44] ^ layer_0[4164]; 
    assign out[1100] = ~(layer_0[3116] ^ layer_0[8540]); 
    assign out[1101] = ~layer_0[5905]; 
    assign out[1102] = ~(layer_0[5217] ^ layer_0[2813]); 
    assign out[1103] = ~layer_0[11408]; 
    assign out[1104] = ~layer_0[23] | (layer_0[23] & layer_0[9296]); 
    assign out[1105] = ~(layer_0[9044] ^ layer_0[8213]); 
    assign out[1106] = layer_0[4780] ^ layer_0[11019]; 
    assign out[1107] = ~(layer_0[8181] ^ layer_0[8475]); 
    assign out[1108] = ~(layer_0[2393] & layer_0[5323]); 
    assign out[1109] = ~(layer_0[8712] ^ layer_0[5944]); 
    assign out[1110] = layer_0[10222] ^ layer_0[9993]; 
    assign out[1111] = layer_0[885] ^ layer_0[11465]; 
    assign out[1112] = layer_0[5514] ^ layer_0[9695]; 
    assign out[1113] = layer_0[5427] | layer_0[11575]; 
    assign out[1114] = layer_0[10846] ^ layer_0[545]; 
    assign out[1115] = layer_0[150] & ~layer_0[9166]; 
    assign out[1116] = layer_0[9598] | layer_0[2797]; 
    assign out[1117] = ~(layer_0[6233] ^ layer_0[6841]); 
    assign out[1118] = ~(layer_0[5364] & layer_0[11237]); 
    assign out[1119] = ~(layer_0[4261] | layer_0[7626]); 
    assign out[1120] = ~layer_0[208]; 
    assign out[1121] = ~(layer_0[387] ^ layer_0[3467]); 
    assign out[1122] = layer_0[2717] ^ layer_0[8927]; 
    assign out[1123] = ~(layer_0[9497] ^ layer_0[1375]); 
    assign out[1124] = layer_0[8112] & ~layer_0[8370]; 
    assign out[1125] = ~(layer_0[5294] ^ layer_0[9910]); 
    assign out[1126] = layer_0[5892] & ~layer_0[9966]; 
    assign out[1127] = ~(layer_0[7665] ^ layer_0[10859]); 
    assign out[1128] = ~layer_0[4833]; 
    assign out[1129] = layer_0[5851] | layer_0[221]; 
    assign out[1130] = ~(layer_0[3007] ^ layer_0[4623]); 
    assign out[1131] = layer_0[4964]; 
    assign out[1132] = ~layer_0[3910]; 
    assign out[1133] = ~(layer_0[9446] | layer_0[3862]); 
    assign out[1134] = layer_0[3769] ^ layer_0[2818]; 
    assign out[1135] = layer_0[9927] & ~layer_0[140]; 
    assign out[1136] = ~(layer_0[3790] ^ layer_0[2864]); 
    assign out[1137] = ~layer_0[10033]; 
    assign out[1138] = layer_0[7823] ^ layer_0[9450]; 
    assign out[1139] = ~layer_0[1597]; 
    assign out[1140] = ~layer_0[756] | (layer_0[756] & layer_0[11065]); 
    assign out[1141] = layer_0[7619] ^ layer_0[1216]; 
    assign out[1142] = layer_0[11058] ^ layer_0[2880]; 
    assign out[1143] = ~layer_0[9627]; 
    assign out[1144] = ~layer_0[672] | (layer_0[672] & layer_0[6326]); 
    assign out[1145] = layer_0[661] & ~layer_0[8385]; 
    assign out[1146] = 1'b0; 
    assign out[1147] = layer_0[4229]; 
    assign out[1148] = ~layer_0[73]; 
    assign out[1149] = ~layer_0[7810] | (layer_0[5511] & layer_0[7810]); 
    assign out[1150] = layer_0[5633] ^ layer_0[9186]; 
    assign out[1151] = ~(layer_0[9966] ^ layer_0[11134]); 
    assign out[1152] = ~(layer_0[2236] ^ layer_0[372]); 
    assign out[1153] = ~(layer_0[5627] ^ layer_0[9850]); 
    assign out[1154] = layer_0[5717]; 
    assign out[1155] = layer_0[2661] | layer_0[5917]; 
    assign out[1156] = ~(layer_0[3674] ^ layer_0[4007]); 
    assign out[1157] = layer_0[10372] & ~layer_0[6710]; 
    assign out[1158] = ~layer_0[5744] | (layer_0[5744] & layer_0[9255]); 
    assign out[1159] = layer_0[9389] ^ layer_0[904]; 
    assign out[1160] = ~(layer_0[7950] & layer_0[845]); 
    assign out[1161] = layer_0[4297] ^ layer_0[3850]; 
    assign out[1162] = ~layer_0[2453]; 
    assign out[1163] = ~(layer_0[3724] ^ layer_0[10818]); 
    assign out[1164] = layer_0[10266]; 
    assign out[1165] = layer_0[10084] & layer_0[6223]; 
    assign out[1166] = layer_0[11194] ^ layer_0[384]; 
    assign out[1167] = ~(layer_0[9200] ^ layer_0[278]); 
    assign out[1168] = ~(layer_0[873] ^ layer_0[9581]); 
    assign out[1169] = layer_0[11653] & ~layer_0[5181]; 
    assign out[1170] = layer_0[227] ^ layer_0[11006]; 
    assign out[1171] = layer_0[11410]; 
    assign out[1172] = layer_0[5687] ^ layer_0[7483]; 
    assign out[1173] = ~layer_0[158]; 
    assign out[1174] = ~(layer_0[10586] ^ layer_0[737]); 
    assign out[1175] = ~(layer_0[4854] ^ layer_0[3026]); 
    assign out[1176] = layer_0[5512]; 
    assign out[1177] = layer_0[8689] & ~layer_0[8543]; 
    assign out[1178] = ~(layer_0[8835] | layer_0[6366]); 
    assign out[1179] = layer_0[5513] ^ layer_0[3923]; 
    assign out[1180] = ~(layer_0[9182] ^ layer_0[5708]); 
    assign out[1181] = layer_0[2615] ^ layer_0[3681]; 
    assign out[1182] = layer_0[2654] ^ layer_0[3638]; 
    assign out[1183] = ~(layer_0[6899] ^ layer_0[9025]); 
    assign out[1184] = ~layer_0[3738]; 
    assign out[1185] = ~(layer_0[1367] ^ layer_0[8316]); 
    assign out[1186] = ~layer_0[874]; 
    assign out[1187] = ~(layer_0[5102] | layer_0[3284]); 
    assign out[1188] = layer_0[11408]; 
    assign out[1189] = layer_0[6341] ^ layer_0[547]; 
    assign out[1190] = ~(layer_0[9958] ^ layer_0[3078]); 
    assign out[1191] = ~layer_0[1293]; 
    assign out[1192] = layer_0[6055] & ~layer_0[11843]; 
    assign out[1193] = layer_0[8446] ^ layer_0[7818]; 
    assign out[1194] = layer_0[4227] ^ layer_0[10239]; 
    assign out[1195] = ~(layer_0[7456] ^ layer_0[7085]); 
    assign out[1196] = ~layer_0[1885]; 
    assign out[1197] = ~(layer_0[11632] & layer_0[8713]); 
    assign out[1198] = layer_0[8183] & layer_0[5334]; 
    assign out[1199] = ~layer_0[994]; 
    assign out[1200] = layer_0[3502]; 
    assign out[1201] = ~(layer_0[4387] ^ layer_0[8719]); 
    assign out[1202] = ~layer_0[6612]; 
    assign out[1203] = layer_0[11730] ^ layer_0[11959]; 
    assign out[1204] = layer_0[5896] & ~layer_0[5292]; 
    assign out[1205] = ~(layer_0[6441] ^ layer_0[1509]); 
    assign out[1206] = layer_0[10535] ^ layer_0[5591]; 
    assign out[1207] = layer_0[5845]; 
    assign out[1208] = ~(layer_0[2120] ^ layer_0[9767]); 
    assign out[1209] = 1'b0; 
    assign out[1210] = layer_0[6928] ^ layer_0[11048]; 
    assign out[1211] = layer_0[7423] & ~layer_0[5035]; 
    assign out[1212] = layer_0[4126] ^ layer_0[7944]; 
    assign out[1213] = ~(layer_0[10878] | layer_0[1829]); 
    assign out[1214] = layer_0[9135] & layer_0[641]; 
    assign out[1215] = ~layer_0[3799] | (layer_0[3799] & layer_0[9857]); 
    assign out[1216] = layer_0[10443] & layer_0[6602]; 
    assign out[1217] = layer_0[3587] & ~layer_0[1816]; 
    assign out[1218] = layer_0[4305] ^ layer_0[10835]; 
    assign out[1219] = layer_0[1864] ^ layer_0[269]; 
    assign out[1220] = layer_0[2392]; 
    assign out[1221] = layer_0[1639] & ~layer_0[3115]; 
    assign out[1222] = layer_0[10346] & layer_0[3110]; 
    assign out[1223] = layer_0[11802] ^ layer_0[9792]; 
    assign out[1224] = ~(layer_0[1031] ^ layer_0[9340]); 
    assign out[1225] = ~(layer_0[4404] ^ layer_0[7243]); 
    assign out[1226] = ~(layer_0[3649] ^ layer_0[9261]); 
    assign out[1227] = layer_0[2335] ^ layer_0[4979]; 
    assign out[1228] = layer_0[4285] & layer_0[8502]; 
    assign out[1229] = layer_0[8515] ^ layer_0[2039]; 
    assign out[1230] = layer_0[10832] | layer_0[2016]; 
    assign out[1231] = layer_0[10244] ^ layer_0[5553]; 
    assign out[1232] = ~layer_0[6239]; 
    assign out[1233] = layer_0[10927] & ~layer_0[8715]; 
    assign out[1234] = layer_0[4975] & layer_0[6800]; 
    assign out[1235] = layer_0[9827]; 
    assign out[1236] = ~layer_0[7201]; 
    assign out[1237] = layer_0[3299] ^ layer_0[2073]; 
    assign out[1238] = layer_0[2928] ^ layer_0[5771]; 
    assign out[1239] = layer_0[8157] ^ layer_0[8167]; 
    assign out[1240] = layer_0[2407] & layer_0[134]; 
    assign out[1241] = ~layer_0[10898] | (layer_0[6916] & layer_0[10898]); 
    assign out[1242] = ~(layer_0[1709] & layer_0[8494]); 
    assign out[1243] = ~(layer_0[4080] ^ layer_0[10063]); 
    assign out[1244] = layer_0[6806]; 
    assign out[1245] = layer_0[3464] & ~layer_0[10120]; 
    assign out[1246] = ~layer_0[1902]; 
    assign out[1247] = layer_0[7485] ^ layer_0[7471]; 
    assign out[1248] = layer_0[6348] & ~layer_0[2783]; 
    assign out[1249] = layer_0[8091] & ~layer_0[11745]; 
    assign out[1250] = ~(layer_0[8517] & layer_0[10413]); 
    assign out[1251] = ~(layer_0[2809] & layer_0[1907]); 
    assign out[1252] = layer_0[1188]; 
    assign out[1253] = ~(layer_0[11662] ^ layer_0[10057]); 
    assign out[1254] = ~(layer_0[3190] ^ layer_0[609]); 
    assign out[1255] = layer_0[271] & ~layer_0[2327]; 
    assign out[1256] = ~(layer_0[4066] | layer_0[6502]); 
    assign out[1257] = layer_0[7361] ^ layer_0[5802]; 
    assign out[1258] = ~layer_0[11151]; 
    assign out[1259] = layer_0[10553] ^ layer_0[11927]; 
    assign out[1260] = ~layer_0[7238] | (layer_0[8796] & layer_0[7238]); 
    assign out[1261] = ~(layer_0[6420] ^ layer_0[4884]); 
    assign out[1262] = layer_0[7875] ^ layer_0[1520]; 
    assign out[1263] = layer_0[8410] ^ layer_0[11052]; 
    assign out[1264] = ~(layer_0[2778] | layer_0[2734]); 
    assign out[1265] = layer_0[6392]; 
    assign out[1266] = layer_0[9737]; 
    assign out[1267] = ~(layer_0[4600] ^ layer_0[2951]); 
    assign out[1268] = ~(layer_0[10845] ^ layer_0[9180]); 
    assign out[1269] = ~(layer_0[11723] ^ layer_0[10374]); 
    assign out[1270] = layer_0[821] & ~layer_0[1344]; 
    assign out[1271] = ~(layer_0[10211] ^ layer_0[2190]); 
    assign out[1272] = ~layer_0[3319]; 
    assign out[1273] = ~layer_0[10795]; 
    assign out[1274] = ~(layer_0[8205] ^ layer_0[1125]); 
    assign out[1275] = layer_0[10737] ^ layer_0[5363]; 
    assign out[1276] = ~(layer_0[11700] & layer_0[2212]); 
    assign out[1277] = ~(layer_0[7821] | layer_0[1349]); 
    assign out[1278] = layer_0[4786] & layer_0[1958]; 
    assign out[1279] = ~layer_0[756]; 
    assign out[1280] = layer_0[2052] & layer_0[10188]; 
    assign out[1281] = layer_0[7655] ^ layer_0[8614]; 
    assign out[1282] = layer_0[8292] ^ layer_0[851]; 
    assign out[1283] = layer_0[5153] & layer_0[993]; 
    assign out[1284] = layer_0[9695] ^ layer_0[5151]; 
    assign out[1285] = layer_0[4163] & ~layer_0[11563]; 
    assign out[1286] = layer_0[10182] & layer_0[346]; 
    assign out[1287] = layer_0[1243] | layer_0[2816]; 
    assign out[1288] = ~(layer_0[2240] ^ layer_0[1227]); 
    assign out[1289] = ~layer_0[10788]; 
    assign out[1290] = layer_0[9272] & layer_0[3586]; 
    assign out[1291] = ~(layer_0[1358] | layer_0[7247]); 
    assign out[1292] = ~(layer_0[4365] ^ layer_0[1542]); 
    assign out[1293] = layer_0[1248] & ~layer_0[479]; 
    assign out[1294] = layer_0[5933] & ~layer_0[350]; 
    assign out[1295] = ~(layer_0[3217] ^ layer_0[4470]); 
    assign out[1296] = layer_0[164] ^ layer_0[10652]; 
    assign out[1297] = ~layer_0[797]; 
    assign out[1298] = ~layer_0[11471] | (layer_0[11471] & layer_0[11200]); 
    assign out[1299] = layer_0[8741] & layer_0[11727]; 
    assign out[1300] = ~(layer_0[2914] ^ layer_0[6506]); 
    assign out[1301] = layer_0[11406] ^ layer_0[1797]; 
    assign out[1302] = layer_0[3864] ^ layer_0[6104]; 
    assign out[1303] = layer_0[468] & ~layer_0[9688]; 
    assign out[1304] = layer_0[11304] ^ layer_0[10656]; 
    assign out[1305] = layer_0[5838] ^ layer_0[8587]; 
    assign out[1306] = ~(layer_0[7075] ^ layer_0[4990]); 
    assign out[1307] = layer_0[789] ^ layer_0[2921]; 
    assign out[1308] = layer_0[8525] ^ layer_0[6281]; 
    assign out[1309] = ~(layer_0[5258] | layer_0[1017]); 
    assign out[1310] = layer_0[8844] & layer_0[330]; 
    assign out[1311] = layer_0[4117]; 
    assign out[1312] = layer_0[8009] | layer_0[5618]; 
    assign out[1313] = ~layer_0[2242]; 
    assign out[1314] = ~layer_0[1337] | (layer_0[1337] & layer_0[4915]); 
    assign out[1315] = ~(layer_0[9626] | layer_0[2144]); 
    assign out[1316] = ~(layer_0[11579] & layer_0[219]); 
    assign out[1317] = layer_0[3782] ^ layer_0[2085]; 
    assign out[1318] = ~(layer_0[1854] ^ layer_0[6566]); 
    assign out[1319] = ~(layer_0[403] ^ layer_0[5129]); 
    assign out[1320] = layer_0[4285] & layer_0[4810]; 
    assign out[1321] = layer_0[3660] ^ layer_0[6149]; 
    assign out[1322] = ~(layer_0[1086] ^ layer_0[11820]); 
    assign out[1323] = ~(layer_0[11794] | layer_0[8444]); 
    assign out[1324] = layer_0[11527]; 
    assign out[1325] = layer_0[3064] ^ layer_0[6183]; 
    assign out[1326] = layer_0[3880] & layer_0[6684]; 
    assign out[1327] = ~layer_0[8343] | (layer_0[8343] & layer_0[10479]); 
    assign out[1328] = layer_0[9983] & ~layer_0[8711]; 
    assign out[1329] = layer_0[9492] ^ layer_0[9776]; 
    assign out[1330] = ~(layer_0[4388] & layer_0[505]); 
    assign out[1331] = ~(layer_0[2192] | layer_0[1293]); 
    assign out[1332] = ~(layer_0[5060] | layer_0[9372]); 
    assign out[1333] = ~layer_0[4870]; 
    assign out[1334] = ~layer_0[6499] | (layer_0[6499] & layer_0[11813]); 
    assign out[1335] = ~(layer_0[1445] ^ layer_0[5346]); 
    assign out[1336] = layer_0[8484]; 
    assign out[1337] = layer_0[7693]; 
    assign out[1338] = layer_0[11079]; 
    assign out[1339] = ~(layer_0[9569] ^ layer_0[1205]); 
    assign out[1340] = ~(layer_0[1671] ^ layer_0[11227]); 
    assign out[1341] = layer_0[4660] ^ layer_0[7558]; 
    assign out[1342] = ~layer_0[7623]; 
    assign out[1343] = ~(layer_0[6517] ^ layer_0[11118]); 
    assign out[1344] = layer_0[8288] & ~layer_0[3041]; 
    assign out[1345] = layer_0[6360] & layer_0[8253]; 
    assign out[1346] = layer_0[6781]; 
    assign out[1347] = layer_0[8383] ^ layer_0[4592]; 
    assign out[1348] = ~layer_0[5261] | (layer_0[5261] & layer_0[1092]); 
    assign out[1349] = ~(layer_0[8038] ^ layer_0[10495]); 
    assign out[1350] = layer_0[8176] & ~layer_0[7258]; 
    assign out[1351] = ~(layer_0[8311] ^ layer_0[8625]); 
    assign out[1352] = ~(layer_0[4777] ^ layer_0[430]); 
    assign out[1353] = ~(layer_0[11177] ^ layer_0[4541]); 
    assign out[1354] = ~layer_0[7211]; 
    assign out[1355] = layer_0[10519] ^ layer_0[6979]; 
    assign out[1356] = layer_0[3869] ^ layer_0[1576]; 
    assign out[1357] = layer_0[8256] & ~layer_0[1764]; 
    assign out[1358] = ~(layer_0[9233] | layer_0[7010]); 
    assign out[1359] = ~(layer_0[3798] ^ layer_0[11862]); 
    assign out[1360] = ~(layer_0[114] ^ layer_0[6063]); 
    assign out[1361] = layer_0[6777] ^ layer_0[11669]; 
    assign out[1362] = ~(layer_0[10293] ^ layer_0[10595]); 
    assign out[1363] = ~(layer_0[3430] ^ layer_0[4552]); 
    assign out[1364] = layer_0[8574] & ~layer_0[5883]; 
    assign out[1365] = ~(layer_0[11292] ^ layer_0[3200]); 
    assign out[1366] = ~(layer_0[4636] & layer_0[7651]); 
    assign out[1367] = layer_0[6597] ^ layer_0[2970]; 
    assign out[1368] = layer_0[10693] ^ layer_0[7206]; 
    assign out[1369] = ~layer_0[6734]; 
    assign out[1370] = ~(layer_0[97] ^ layer_0[8848]); 
    assign out[1371] = layer_0[5837] ^ layer_0[2340]; 
    assign out[1372] = ~(layer_0[6591] | layer_0[3706]); 
    assign out[1373] = layer_0[5544]; 
    assign out[1374] = ~layer_0[4284]; 
    assign out[1375] = layer_0[517] & ~layer_0[3112]; 
    assign out[1376] = layer_0[3888] & ~layer_0[9061]; 
    assign out[1377] = ~layer_0[2421]; 
    assign out[1378] = layer_0[8260] & layer_0[11776]; 
    assign out[1379] = ~layer_0[4469]; 
    assign out[1380] = ~layer_0[10521]; 
    assign out[1381] = layer_0[11509] ^ layer_0[3636]; 
    assign out[1382] = ~(layer_0[486] ^ layer_0[4967]); 
    assign out[1383] = layer_0[2571] & layer_0[733]; 
    assign out[1384] = ~layer_0[1281]; 
    assign out[1385] = ~layer_0[2012] | (layer_0[2823] & layer_0[2012]); 
    assign out[1386] = ~layer_0[11625] | (layer_0[11625] & layer_0[6866]); 
    assign out[1387] = ~layer_0[82] | (layer_0[8023] & layer_0[82]); 
    assign out[1388] = layer_0[5616] ^ layer_0[9576]; 
    assign out[1389] = layer_0[11004] ^ layer_0[2917]; 
    assign out[1390] = ~layer_0[8851]; 
    assign out[1391] = ~layer_0[6609]; 
    assign out[1392] = layer_0[4747]; 
    assign out[1393] = ~(layer_0[3585] ^ layer_0[9932]); 
    assign out[1394] = ~(layer_0[4580] ^ layer_0[3651]); 
    assign out[1395] = layer_0[4956] & ~layer_0[7984]; 
    assign out[1396] = ~(layer_0[3938] | layer_0[1723]); 
    assign out[1397] = ~(layer_0[8148] ^ layer_0[11560]); 
    assign out[1398] = layer_0[294] ^ layer_0[2996]; 
    assign out[1399] = ~(layer_0[153] ^ layer_0[7047]); 
    assign out[1400] = layer_0[4374] ^ layer_0[10688]; 
    assign out[1401] = ~layer_0[1103]; 
    assign out[1402] = ~(layer_0[9722] ^ layer_0[4976]); 
    assign out[1403] = layer_0[11303] ^ layer_0[6225]; 
    assign out[1404] = ~layer_0[2801]; 
    assign out[1405] = layer_0[9156] ^ layer_0[2979]; 
    assign out[1406] = ~(layer_0[2074] ^ layer_0[4563]); 
    assign out[1407] = ~(layer_0[10029] ^ layer_0[11919]); 
    assign out[1408] = layer_0[1468] ^ layer_0[5091]; 
    assign out[1409] = ~(layer_0[3018] & layer_0[9541]); 
    assign out[1410] = layer_0[10765] & layer_0[5855]; 
    assign out[1411] = ~layer_0[3442]; 
    assign out[1412] = layer_0[1583]; 
    assign out[1413] = ~(layer_0[7193] ^ layer_0[8827]); 
    assign out[1414] = layer_0[3697] & ~layer_0[11024]; 
    assign out[1415] = ~(layer_0[3715] ^ layer_0[3644]); 
    assign out[1416] = layer_0[7962] ^ layer_0[568]; 
    assign out[1417] = layer_0[8293] ^ layer_0[7914]; 
    assign out[1418] = layer_0[11552] ^ layer_0[10222]; 
    assign out[1419] = ~layer_0[10153]; 
    assign out[1420] = ~layer_0[6634]; 
    assign out[1421] = ~(layer_0[6844] ^ layer_0[2307]); 
    assign out[1422] = ~layer_0[3682]; 
    assign out[1423] = layer_0[8897] & ~layer_0[7268]; 
    assign out[1424] = layer_0[7224] ^ layer_0[5590]; 
    assign out[1425] = layer_0[7174] ^ layer_0[3686]; 
    assign out[1426] = layer_0[10641] & ~layer_0[11936]; 
    assign out[1427] = ~(layer_0[4900] ^ layer_0[6265]); 
    assign out[1428] = layer_0[1428] ^ layer_0[9759]; 
    assign out[1429] = layer_0[6980] & ~layer_0[3695]; 
    assign out[1430] = layer_0[2441] ^ layer_0[2955]; 
    assign out[1431] = ~(layer_0[6614] ^ layer_0[10338]); 
    assign out[1432] = layer_0[2423] & ~layer_0[1156]; 
    assign out[1433] = layer_0[9053] ^ layer_0[6681]; 
    assign out[1434] = layer_0[4345] ^ layer_0[7631]; 
    assign out[1435] = ~(layer_0[5980] | layer_0[10160]); 
    assign out[1436] = ~layer_0[3160]; 
    assign out[1437] = ~layer_0[9872]; 
    assign out[1438] = layer_0[9154] ^ layer_0[9726]; 
    assign out[1439] = layer_0[3607] ^ layer_0[4522]; 
    assign out[1440] = ~(layer_0[2417] ^ layer_0[7174]); 
    assign out[1441] = layer_0[9032]; 
    assign out[1442] = ~(layer_0[7592] | layer_0[7696]); 
    assign out[1443] = ~layer_0[9691]; 
    assign out[1444] = layer_0[4809] ^ layer_0[7873]; 
    assign out[1445] = layer_0[9959] ^ layer_0[7859]; 
    assign out[1446] = ~(layer_0[6660] ^ layer_0[5301]); 
    assign out[1447] = layer_0[6693] ^ layer_0[1476]; 
    assign out[1448] = ~(layer_0[6017] ^ layer_0[2931]); 
    assign out[1449] = layer_0[3149]; 
    assign out[1450] = layer_0[6961]; 
    assign out[1451] = ~(layer_0[5798] ^ layer_0[3629]); 
    assign out[1452] = layer_0[11404] ^ layer_0[4662]; 
    assign out[1453] = layer_0[10884] ^ layer_0[1373]; 
    assign out[1454] = layer_0[7620] & ~layer_0[9092]; 
    assign out[1455] = ~layer_0[11290] | (layer_0[11290] & layer_0[7463]); 
    assign out[1456] = ~(layer_0[1005] ^ layer_0[7473]); 
    assign out[1457] = ~(layer_0[6915] ^ layer_0[1782]); 
    assign out[1458] = layer_0[1128]; 
    assign out[1459] = layer_0[11162] & ~layer_0[8042]; 
    assign out[1460] = ~layer_0[9369] | (layer_0[9369] & layer_0[1319]); 
    assign out[1461] = ~(layer_0[7980] ^ layer_0[10340]); 
    assign out[1462] = ~layer_0[73] | (layer_0[6374] & layer_0[73]); 
    assign out[1463] = ~(layer_0[10783] ^ layer_0[10643]); 
    assign out[1464] = ~(layer_0[6037] ^ layer_0[3359]); 
    assign out[1465] = ~(layer_0[2167] ^ layer_0[573]); 
    assign out[1466] = layer_0[10702]; 
    assign out[1467] = layer_0[1088] & ~layer_0[3992]; 
    assign out[1468] = layer_0[6494] ^ layer_0[10813]; 
    assign out[1469] = layer_0[8504] ^ layer_0[945]; 
    assign out[1470] = layer_0[8884] ^ layer_0[1587]; 
    assign out[1471] = layer_0[6250] & ~layer_0[7768]; 
    assign out[1472] = ~(layer_0[2456] | layer_0[10359]); 
    assign out[1473] = layer_0[5032]; 
    assign out[1474] = ~(layer_0[10642] | layer_0[6745]); 
    assign out[1475] = ~layer_0[10660]; 
    assign out[1476] = ~layer_0[2157]; 
    assign out[1477] = layer_0[6246]; 
    assign out[1478] = layer_0[2513] & ~layer_0[4204]; 
    assign out[1479] = ~(layer_0[7557] ^ layer_0[8654]); 
    assign out[1480] = layer_0[11480] & ~layer_0[759]; 
    assign out[1481] = ~(layer_0[6579] ^ layer_0[2369]); 
    assign out[1482] = layer_0[7544]; 
    assign out[1483] = ~layer_0[7450] | (layer_0[7450] & layer_0[8050]); 
    assign out[1484] = ~layer_0[2448]; 
    assign out[1485] = ~(layer_0[3072] | layer_0[10367]); 
    assign out[1486] = layer_0[4423]; 
    assign out[1487] = layer_0[8907] ^ layer_0[11829]; 
    assign out[1488] = layer_0[3088]; 
    assign out[1489] = layer_0[1444] & ~layer_0[2627]; 
    assign out[1490] = ~(layer_0[9444] ^ layer_0[411]); 
    assign out[1491] = layer_0[429] ^ layer_0[3630]; 
    assign out[1492] = layer_0[1011] & ~layer_0[3664]; 
    assign out[1493] = ~layer_0[3667]; 
    assign out[1494] = ~layer_0[11353] | (layer_0[11353] & layer_0[8709]); 
    assign out[1495] = ~layer_0[5503]; 
    assign out[1496] = layer_0[5083] & layer_0[1271]; 
    assign out[1497] = ~layer_0[4921]; 
    assign out[1498] = layer_0[513] & ~layer_0[11053]; 
    assign out[1499] = ~layer_0[9664] | (layer_0[9664] & layer_0[4535]); 
    assign out[1500] = layer_0[3094] & ~layer_0[1399]; 
    assign out[1501] = ~(layer_0[6029] ^ layer_0[6713]); 
    assign out[1502] = ~(layer_0[9208] ^ layer_0[3027]); 
    assign out[1503] = layer_0[2904]; 
    assign out[1504] = layer_0[2642] ^ layer_0[8510]; 
    assign out[1505] = ~(layer_0[8014] ^ layer_0[7386]); 
    assign out[1506] = layer_0[6736]; 
    assign out[1507] = ~layer_0[6516]; 
    assign out[1508] = layer_0[7687] ^ layer_0[256]; 
    assign out[1509] = layer_0[1260]; 
    assign out[1510] = layer_0[7420] ^ layer_0[9481]; 
    assign out[1511] = layer_0[8831] ^ layer_0[2095]; 
    assign out[1512] = ~(layer_0[4135] ^ layer_0[10432]); 
    assign out[1513] = layer_0[1443] ^ layer_0[946]; 
    assign out[1514] = layer_0[9031] | layer_0[11189]; 
    assign out[1515] = ~(layer_0[11901] | layer_0[5141]); 
    assign out[1516] = ~(layer_0[1087] ^ layer_0[9560]); 
    assign out[1517] = ~layer_0[7955]; 
    assign out[1518] = ~layer_0[9815]; 
    assign out[1519] = layer_0[5589] & ~layer_0[10217]; 
    assign out[1520] = ~(layer_0[4628] | layer_0[9136]); 
    assign out[1521] = layer_0[6505] ^ layer_0[10540]; 
    assign out[1522] = layer_0[7266] ^ layer_0[8635]; 
    assign out[1523] = ~(layer_0[4929] ^ layer_0[3187]); 
    assign out[1524] = layer_0[6548]; 
    assign out[1525] = ~(layer_0[1051] ^ layer_0[10176]); 
    assign out[1526] = ~layer_0[4544]; 
    assign out[1527] = ~(layer_0[1936] ^ layer_0[5097]); 
    assign out[1528] = ~(layer_0[8663] | layer_0[8051]); 
    assign out[1529] = ~(layer_0[8878] & layer_0[11533]); 
    assign out[1530] = ~(layer_0[4182] ^ layer_0[11470]); 
    assign out[1531] = ~(layer_0[3053] | layer_0[1197]); 
    assign out[1532] = ~(layer_0[7809] ^ layer_0[695]); 
    assign out[1533] = layer_0[4863]; 
    assign out[1534] = layer_0[6144] & layer_0[5189]; 
    assign out[1535] = layer_0[11881] ^ layer_0[7411]; 
    assign out[1536] = ~(layer_0[3304] ^ layer_0[2545]); 
    assign out[1537] = ~(layer_0[9731] ^ layer_0[1990]); 
    assign out[1538] = layer_0[5401]; 
    assign out[1539] = layer_0[9137] & ~layer_0[4639]; 
    assign out[1540] = layer_0[6063]; 
    assign out[1541] = ~layer_0[5373]; 
    assign out[1542] = ~(layer_0[9259] ^ layer_0[6816]); 
    assign out[1543] = layer_0[562]; 
    assign out[1544] = layer_0[1378] ^ layer_0[8922]; 
    assign out[1545] = layer_0[1193] ^ layer_0[8405]; 
    assign out[1546] = ~(layer_0[2987] ^ layer_0[1319]); 
    assign out[1547] = ~(layer_0[5086] ^ layer_0[2478]); 
    assign out[1548] = ~(layer_0[2796] & layer_0[6536]); 
    assign out[1549] = ~(layer_0[4133] ^ layer_0[3247]); 
    assign out[1550] = layer_0[10128] & ~layer_0[4416]; 
    assign out[1551] = ~(layer_0[2969] | layer_0[3895]); 
    assign out[1552] = layer_0[163]; 
    assign out[1553] = ~(layer_0[10231] ^ layer_0[5541]); 
    assign out[1554] = ~(layer_0[9681] | layer_0[3872]); 
    assign out[1555] = layer_0[9969] ^ layer_0[5363]; 
    assign out[1556] = ~(layer_0[9682] ^ layer_0[4894]); 
    assign out[1557] = layer_0[7049] & layer_0[5976]; 
    assign out[1558] = ~(layer_0[11226] ^ layer_0[9354]); 
    assign out[1559] = ~(layer_0[5229] & layer_0[11963]); 
    assign out[1560] = layer_0[4062] ^ layer_0[10551]; 
    assign out[1561] = ~layer_0[3248] | (layer_0[3248] & layer_0[9418]); 
    assign out[1562] = layer_0[10137] ^ layer_0[6821]; 
    assign out[1563] = ~(layer_0[7402] ^ layer_0[5107]); 
    assign out[1564] = ~(layer_0[9125] ^ layer_0[7133]); 
    assign out[1565] = ~(layer_0[6054] ^ layer_0[4597]); 
    assign out[1566] = ~layer_0[10030] | (layer_0[3558] & layer_0[10030]); 
    assign out[1567] = layer_0[619] ^ layer_0[7507]; 
    assign out[1568] = ~(layer_0[548] | layer_0[4390]); 
    assign out[1569] = layer_0[2491]; 
    assign out[1570] = ~(layer_0[10780] ^ layer_0[3638]); 
    assign out[1571] = ~(layer_0[11915] | layer_0[1551]); 
    assign out[1572] = layer_0[11529] ^ layer_0[3631]; 
    assign out[1573] = layer_0[8433] & ~layer_0[806]; 
    assign out[1574] = layer_0[7505] & layer_0[4748]; 
    assign out[1575] = ~layer_0[10824]; 
    assign out[1576] = ~(layer_0[2028] ^ layer_0[2019]); 
    assign out[1577] = layer_0[4056] & ~layer_0[8147]; 
    assign out[1578] = layer_0[10632] ^ layer_0[3541]; 
    assign out[1579] = layer_0[11605] ^ layer_0[8608]; 
    assign out[1580] = layer_0[7777] ^ layer_0[9599]; 
    assign out[1581] = layer_0[11618] | layer_0[5923]; 
    assign out[1582] = ~layer_0[4789]; 
    assign out[1583] = layer_0[7644] ^ layer_0[3099]; 
    assign out[1584] = ~layer_0[4665]; 
    assign out[1585] = ~(layer_0[3038] ^ layer_0[10700]); 
    assign out[1586] = layer_0[4436] ^ layer_0[4399]; 
    assign out[1587] = ~layer_0[162]; 
    assign out[1588] = ~(layer_0[3321] ^ layer_0[10451]); 
    assign out[1589] = ~layer_0[10304]; 
    assign out[1590] = ~(layer_0[3490] ^ layer_0[11694]); 
    assign out[1591] = ~layer_0[10681]; 
    assign out[1592] = ~layer_0[4989]; 
    assign out[1593] = ~layer_0[8428]; 
    assign out[1594] = ~(layer_0[9696] ^ layer_0[3617]); 
    assign out[1595] = layer_0[8988] ^ layer_0[9781]; 
    assign out[1596] = ~(layer_0[3709] ^ layer_0[56]); 
    assign out[1597] = layer_0[11354]; 
    assign out[1598] = layer_0[637] ^ layer_0[10105]; 
    assign out[1599] = layer_0[2755] & ~layer_0[8067]; 
    assign out[1600] = ~(layer_0[9885] ^ layer_0[4464]); 
    assign out[1601] = layer_0[3878]; 
    assign out[1602] = ~(layer_0[4166] ^ layer_0[9956]); 
    assign out[1603] = layer_0[761] ^ layer_0[10333]; 
    assign out[1604] = ~(layer_0[449] ^ layer_0[3671]); 
    assign out[1605] = ~(layer_0[6836] ^ layer_0[8509]); 
    assign out[1606] = ~(layer_0[1759] ^ layer_0[8372]); 
    assign out[1607] = ~(layer_0[3029] ^ layer_0[7699]); 
    assign out[1608] = ~layer_0[1857]; 
    assign out[1609] = layer_0[8607] ^ layer_0[3972]; 
    assign out[1610] = ~(layer_0[7627] | layer_0[11910]); 
    assign out[1611] = layer_0[9036] & ~layer_0[11234]; 
    assign out[1612] = ~(layer_0[3046] | layer_0[3251]); 
    assign out[1613] = ~layer_0[1312] | (layer_0[1312] & layer_0[1194]); 
    assign out[1614] = ~(layer_0[5500] ^ layer_0[10575]); 
    assign out[1615] = ~layer_0[5834]; 
    assign out[1616] = ~layer_0[5358] | (layer_0[830] & layer_0[5358]); 
    assign out[1617] = ~layer_0[1698]; 
    assign out[1618] = ~(layer_0[9825] ^ layer_0[7845]); 
    assign out[1619] = ~(layer_0[4940] | layer_0[8409]); 
    assign out[1620] = ~layer_0[1420]; 
    assign out[1621] = layer_0[8226]; 
    assign out[1622] = layer_0[2092] ^ layer_0[5075]; 
    assign out[1623] = layer_0[11091] | layer_0[6886]; 
    assign out[1624] = ~(layer_0[10947] ^ layer_0[9773]); 
    assign out[1625] = ~(layer_0[1693] | layer_0[10228]); 
    assign out[1626] = ~(layer_0[2958] ^ layer_0[7171]); 
    assign out[1627] = ~layer_0[308]; 
    assign out[1628] = layer_0[5458] ^ layer_0[4347]; 
    assign out[1629] = layer_0[1300]; 
    assign out[1630] = layer_0[7441] & ~layer_0[9918]; 
    assign out[1631] = layer_0[8942] & ~layer_0[2879]; 
    assign out[1632] = layer_0[3520] & ~layer_0[5340]; 
    assign out[1633] = layer_0[6446] ^ layer_0[7058]; 
    assign out[1634] = ~(layer_0[5038] | layer_0[8568]); 
    assign out[1635] = ~layer_0[198]; 
    assign out[1636] = layer_0[8811] ^ layer_0[4064]; 
    assign out[1637] = layer_0[5148] | layer_0[2383]; 
    assign out[1638] = ~layer_0[3283] | (layer_0[3283] & layer_0[1593]); 
    assign out[1639] = layer_0[550]; 
    assign out[1640] = layer_0[989] ^ layer_0[2709]; 
    assign out[1641] = layer_0[7044] ^ layer_0[9559]; 
    assign out[1642] = ~layer_0[6955] | (layer_0[6955] & layer_0[2820]); 
    assign out[1643] = layer_0[7303] ^ layer_0[2596]; 
    assign out[1644] = ~(layer_0[898] | layer_0[940]); 
    assign out[1645] = ~(layer_0[1200] ^ layer_0[6620]); 
    assign out[1646] = ~layer_0[8798] | (layer_0[9064] & layer_0[8798]); 
    assign out[1647] = ~(layer_0[1038] ^ layer_0[4434]); 
    assign out[1648] = ~(layer_0[1754] ^ layer_0[10786]); 
    assign out[1649] = ~(layer_0[11214] | layer_0[1240]); 
    assign out[1650] = layer_0[7904] ^ layer_0[7442]; 
    assign out[1651] = ~layer_0[11064]; 
    assign out[1652] = layer_0[6373]; 
    assign out[1653] = layer_0[270] & ~layer_0[1794]; 
    assign out[1654] = layer_0[4200] ^ layer_0[7143]; 
    assign out[1655] = ~(layer_0[9074] ^ layer_0[3867]); 
    assign out[1656] = layer_0[4229] & layer_0[8895]; 
    assign out[1657] = ~layer_0[1696]; 
    assign out[1658] = ~(layer_0[1811] ^ layer_0[7776]); 
    assign out[1659] = layer_0[9926]; 
    assign out[1660] = layer_0[5739] & ~layer_0[9851]; 
    assign out[1661] = layer_0[8552]; 
    assign out[1662] = layer_0[8577] & ~layer_0[1759]; 
    assign out[1663] = ~(layer_0[3410] ^ layer_0[5938]); 
    assign out[1664] = layer_0[8319]; 
    assign out[1665] = ~(layer_0[4422] ^ layer_0[6452]); 
    assign out[1666] = layer_0[3954] ^ layer_0[4299]; 
    assign out[1667] = layer_0[3800] & ~layer_0[5001]; 
    assign out[1668] = layer_0[10447] ^ layer_0[4189]; 
    assign out[1669] = layer_0[3760] ^ layer_0[5227]; 
    assign out[1670] = ~layer_0[11032]; 
    assign out[1671] = layer_0[1626] ^ layer_0[8641]; 
    assign out[1672] = layer_0[5368] ^ layer_0[11093]; 
    assign out[1673] = layer_0[2230] ^ layer_0[10194]; 
    assign out[1674] = layer_0[635]; 
    assign out[1675] = ~(layer_0[9606] ^ layer_0[1248]); 
    assign out[1676] = layer_0[2283]; 
    assign out[1677] = ~layer_0[3831]; 
    assign out[1678] = ~(layer_0[2119] ^ layer_0[3464]); 
    assign out[1679] = ~(layer_0[2973] ^ layer_0[2713]); 
    assign out[1680] = layer_0[5603] ^ layer_0[4701]; 
    assign out[1681] = layer_0[614] & ~layer_0[7262]; 
    assign out[1682] = layer_0[5586] & layer_0[10993]; 
    assign out[1683] = ~(layer_0[5121] ^ layer_0[1311]); 
    assign out[1684] = ~(layer_0[118] ^ layer_0[5215]); 
    assign out[1685] = layer_0[11606]; 
    assign out[1686] = ~(layer_0[6019] ^ layer_0[8683]); 
    assign out[1687] = layer_0[7592] ^ layer_0[5791]; 
    assign out[1688] = layer_0[8599] ^ layer_0[10766]; 
    assign out[1689] = ~(layer_0[5223] ^ layer_0[8610]); 
    assign out[1690] = layer_0[5172] ^ layer_0[608]; 
    assign out[1691] = layer_0[464] ^ layer_0[1621]; 
    assign out[1692] = ~(layer_0[1650] ^ layer_0[9037]); 
    assign out[1693] = layer_0[4087] ^ layer_0[3998]; 
    assign out[1694] = ~(layer_0[7381] ^ layer_0[8579]); 
    assign out[1695] = layer_0[7281] & ~layer_0[5392]; 
    assign out[1696] = layer_0[4608] ^ layer_0[4508]; 
    assign out[1697] = ~(layer_0[11812] & layer_0[359]); 
    assign out[1698] = layer_0[4129] & layer_0[7167]; 
    assign out[1699] = layer_0[656] & ~layer_0[5724]; 
    assign out[1700] = layer_0[7064] & ~layer_0[5825]; 
    assign out[1701] = layer_0[4775] ^ layer_0[3658]; 
    assign out[1702] = ~(layer_0[10223] ^ layer_0[1818]); 
    assign out[1703] = layer_0[4852] ^ layer_0[4670]; 
    assign out[1704] = layer_0[4275] ^ layer_0[8613]; 
    assign out[1705] = ~layer_0[6116] | (layer_0[273] & layer_0[6116]); 
    assign out[1706] = layer_0[5601] ^ layer_0[2383]; 
    assign out[1707] = ~(layer_0[5367] ^ layer_0[10684]); 
    assign out[1708] = layer_0[10491] ^ layer_0[5222]; 
    assign out[1709] = layer_0[10636] & ~layer_0[8655]; 
    assign out[1710] = layer_0[7376]; 
    assign out[1711] = ~(layer_0[5844] ^ layer_0[1120]); 
    assign out[1712] = ~(layer_0[11960] ^ layer_0[3212]); 
    assign out[1713] = ~(layer_0[991] & layer_0[7757]); 
    assign out[1714] = layer_0[3701] ^ layer_0[6972]; 
    assign out[1715] = layer_0[1677] ^ layer_0[10755]; 
    assign out[1716] = ~(layer_0[1604] ^ layer_0[2957]); 
    assign out[1717] = ~layer_0[8596]; 
    assign out[1718] = ~(layer_0[8985] ^ layer_0[9703]); 
    assign out[1719] = ~(layer_0[8547] | layer_0[10023]); 
    assign out[1720] = ~(layer_0[9343] ^ layer_0[3871]); 
    assign out[1721] = layer_0[786] & ~layer_0[5069]; 
    assign out[1722] = layer_0[8064] & layer_0[8312]; 
    assign out[1723] = layer_0[1850] ^ layer_0[2776]; 
    assign out[1724] = ~(layer_0[10543] ^ layer_0[5026]); 
    assign out[1725] = ~(layer_0[11020] ^ layer_0[3659]); 
    assign out[1726] = layer_0[3658] ^ layer_0[3086]; 
    assign out[1727] = layer_0[5165] ^ layer_0[11121]; 
    assign out[1728] = layer_0[601] ^ layer_0[4286]; 
    assign out[1729] = layer_0[11109] & layer_0[6682]; 
    assign out[1730] = ~(layer_0[11978] ^ layer_0[7846]); 
    assign out[1731] = layer_0[8643] ^ layer_0[605]; 
    assign out[1732] = ~(layer_0[11057] | layer_0[7819]); 
    assign out[1733] = layer_0[8015]; 
    assign out[1734] = ~(layer_0[10619] | layer_0[7958]); 
    assign out[1735] = layer_0[6938] ^ layer_0[11590]; 
    assign out[1736] = ~(layer_0[5637] ^ layer_0[8560]); 
    assign out[1737] = ~(layer_0[1486] ^ layer_0[8846]); 
    assign out[1738] = ~(layer_0[2856] ^ layer_0[7057]); 
    assign out[1739] = ~(layer_0[1366] ^ layer_0[6087]); 
    assign out[1740] = ~(layer_0[1743] ^ layer_0[3733]); 
    assign out[1741] = ~(layer_0[5341] ^ layer_0[8007]); 
    assign out[1742] = layer_0[11254] ^ layer_0[10531]; 
    assign out[1743] = ~(layer_0[3834] ^ layer_0[2187]); 
    assign out[1744] = layer_0[9127] ^ layer_0[11111]; 
    assign out[1745] = ~(layer_0[7099] | layer_0[1302]); 
    assign out[1746] = ~(layer_0[10685] ^ layer_0[3584]); 
    assign out[1747] = layer_0[4013] ^ layer_0[6498]; 
    assign out[1748] = ~(layer_0[7944] ^ layer_0[11635]); 
    assign out[1749] = ~(layer_0[6973] ^ layer_0[3364]); 
    assign out[1750] = ~(layer_0[7114] ^ layer_0[613]); 
    assign out[1751] = ~(layer_0[5641] ^ layer_0[9669]); 
    assign out[1752] = layer_0[2100] ^ layer_0[7702]; 
    assign out[1753] = layer_0[3885] ^ layer_0[6549]; 
    assign out[1754] = ~(layer_0[8861] ^ layer_0[2043]); 
    assign out[1755] = ~layer_0[11481]; 
    assign out[1756] = layer_0[10041] ^ layer_0[8979]; 
    assign out[1757] = ~(layer_0[3243] ^ layer_0[5916]); 
    assign out[1758] = ~(layer_0[4362] ^ layer_0[2740]); 
    assign out[1759] = ~(layer_0[11987] ^ layer_0[3955]); 
    assign out[1760] = ~(layer_0[4468] | layer_0[1092]); 
    assign out[1761] = layer_0[2867] & ~layer_0[8309]; 
    assign out[1762] = ~(layer_0[10100] ^ layer_0[5269]); 
    assign out[1763] = layer_0[1630] ^ layer_0[3437]; 
    assign out[1764] = layer_0[4977] & layer_0[10068]; 
    assign out[1765] = ~(layer_0[10612] | layer_0[11812]); 
    assign out[1766] = layer_0[2379] ^ layer_0[11776]; 
    assign out[1767] = ~(layer_0[7982] ^ layer_0[8745]); 
    assign out[1768] = ~layer_0[951] | (layer_0[951] & layer_0[5238]); 
    assign out[1769] = layer_0[2246] & layer_0[10767]; 
    assign out[1770] = ~(layer_0[4558] ^ layer_0[5202]); 
    assign out[1771] = ~(layer_0[648] ^ layer_0[10051]); 
    assign out[1772] = ~(layer_0[11230] | layer_0[11908]); 
    assign out[1773] = ~(layer_0[3456] & layer_0[9923]); 
    assign out[1774] = layer_0[7361] ^ layer_0[293]; 
    assign out[1775] = layer_0[10566]; 
    assign out[1776] = ~layer_0[5524] | (layer_0[5524] & layer_0[8645]); 
    assign out[1777] = ~layer_0[7676]; 
    assign out[1778] = layer_0[11858] ^ layer_0[10469]; 
    assign out[1779] = layer_0[872] ^ layer_0[9911]; 
    assign out[1780] = layer_0[8678]; 
    assign out[1781] = ~(layer_0[7357] ^ layer_0[2071]); 
    assign out[1782] = layer_0[2753]; 
    assign out[1783] = layer_0[10650] & layer_0[10802]; 
    assign out[1784] = ~(layer_0[9081] ^ layer_0[8599]); 
    assign out[1785] = ~layer_0[10824]; 
    assign out[1786] = ~(layer_0[10678] ^ layer_0[10235]); 
    assign out[1787] = layer_0[3892] ^ layer_0[4015]; 
    assign out[1788] = layer_0[1731] ^ layer_0[11440]; 
    assign out[1789] = layer_0[4611]; 
    assign out[1790] = layer_0[209] & ~layer_0[1963]; 
    assign out[1791] = layer_0[10881] & ~layer_0[441]; 
    assign out[1792] = ~layer_0[3375]; 
    assign out[1793] = layer_0[9506] ^ layer_0[1362]; 
    assign out[1794] = layer_0[4528] ^ layer_0[9630]; 
    assign out[1795] = layer_0[9128] ^ layer_0[2610]; 
    assign out[1796] = ~layer_0[2390]; 
    assign out[1797] = ~(layer_0[4621] | layer_0[6921]); 
    assign out[1798] = ~layer_0[5311] | (layer_0[11671] & layer_0[5311]); 
    assign out[1799] = layer_0[8785] | layer_0[2335]; 
    assign out[1800] = ~(layer_0[8883] ^ layer_0[5863]); 
    assign out[1801] = ~(layer_0[10108] ^ layer_0[9311]); 
    assign out[1802] = layer_0[7932] ^ layer_0[620]; 
    assign out[1803] = layer_0[10408] & ~layer_0[1735]; 
    assign out[1804] = ~layer_0[1460]; 
    assign out[1805] = ~(layer_0[10580] ^ layer_0[10135]); 
    assign out[1806] = ~(layer_0[10157] ^ layer_0[6075]); 
    assign out[1807] = ~(layer_0[11864] ^ layer_0[6287]); 
    assign out[1808] = ~(layer_0[2048] ^ layer_0[10287]); 
    assign out[1809] = ~(layer_0[2262] ^ layer_0[7688]); 
    assign out[1810] = layer_0[10259] & layer_0[7350]; 
    assign out[1811] = layer_0[10358] ^ layer_0[8032]; 
    assign out[1812] = ~layer_0[10462]; 
    assign out[1813] = ~(layer_0[153] ^ layer_0[8000]); 
    assign out[1814] = layer_0[3125] & ~layer_0[3915]; 
    assign out[1815] = ~(layer_0[8799] ^ layer_0[6001]); 
    assign out[1816] = layer_0[4192] ^ layer_0[10066]; 
    assign out[1817] = layer_0[4444] ^ layer_0[4675]; 
    assign out[1818] = 1'b0; 
    assign out[1819] = layer_0[4843] ^ layer_0[5974]; 
    assign out[1820] = layer_0[9687] ^ layer_0[7658]; 
    assign out[1821] = ~(layer_0[7341] ^ layer_0[8369]); 
    assign out[1822] = ~layer_0[9543]; 
    assign out[1823] = ~(layer_0[1347] ^ layer_0[6153]); 
    assign out[1824] = ~(layer_0[1261] | layer_0[11854]); 
    assign out[1825] = ~layer_0[1340] | (layer_0[1340] & layer_0[7325]); 
    assign out[1826] = layer_0[2329] | layer_0[9803]; 
    assign out[1827] = ~(layer_0[1455] ^ layer_0[1801]); 
    assign out[1828] = layer_0[11655] & layer_0[2828]; 
    assign out[1829] = layer_0[98] & ~layer_0[11230]; 
    assign out[1830] = layer_0[8295] ^ layer_0[6913]; 
    assign out[1831] = ~(layer_0[6390] ^ layer_0[5609]); 
    assign out[1832] = ~(layer_0[3016] ^ layer_0[10690]); 
    assign out[1833] = layer_0[4426] | layer_0[861]; 
    assign out[1834] = layer_0[4855]; 
    assign out[1835] = layer_0[2986] & ~layer_0[2464]; 
    assign out[1836] = layer_0[7253] & ~layer_0[10228]; 
    assign out[1837] = ~(layer_0[2999] ^ layer_0[4558]); 
    assign out[1838] = ~layer_0[11804]; 
    assign out[1839] = layer_0[5155] & ~layer_0[8247]; 
    assign out[1840] = layer_0[1228] & ~layer_0[4400]; 
    assign out[1841] = ~(layer_0[4457] ^ layer_0[6616]); 
    assign out[1842] = layer_0[5396] ^ layer_0[4063]; 
    assign out[1843] = ~(layer_0[10362] ^ layer_0[9739]); 
    assign out[1844] = layer_0[7022] ^ layer_0[8878]; 
    assign out[1845] = layer_0[10230] & layer_0[1701]; 
    assign out[1846] = layer_0[1564] & ~layer_0[267]; 
    assign out[1847] = ~layer_0[3951]; 
    assign out[1848] = ~(layer_0[840] ^ layer_0[11638]); 
    assign out[1849] = layer_0[2361] & ~layer_0[3164]; 
    assign out[1850] = ~(layer_0[8239] ^ layer_0[2054]); 
    assign out[1851] = ~(layer_0[10633] | layer_0[7462]); 
    assign out[1852] = layer_0[7053] & ~layer_0[5830]; 
    assign out[1853] = ~(layer_0[5188] ^ layer_0[8300]); 
    assign out[1854] = ~(layer_0[9062] ^ layer_0[4806]); 
    assign out[1855] = layer_0[10969] ^ layer_0[5732]; 
    assign out[1856] = ~(layer_0[5015] | layer_0[11403]); 
    assign out[1857] = ~(layer_0[3764] ^ layer_0[8665]); 
    assign out[1858] = layer_0[2812] ^ layer_0[7221]; 
    assign out[1859] = layer_0[5887] | layer_0[11846]; 
    assign out[1860] = layer_0[916] & ~layer_0[7756]; 
    assign out[1861] = layer_0[7230] & ~layer_0[8177]; 
    assign out[1862] = layer_0[11251] ^ layer_0[5947]; 
    assign out[1863] = layer_0[8945] ^ layer_0[7523]; 
    assign out[1864] = layer_0[11993] ^ layer_0[5025]; 
    assign out[1865] = ~(layer_0[10201] ^ layer_0[7941]); 
    assign out[1866] = layer_0[9001] ^ layer_0[2388]; 
    assign out[1867] = ~(layer_0[9960] & layer_0[8214]); 
    assign out[1868] = ~(layer_0[9185] ^ layer_0[1866]); 
    assign out[1869] = layer_0[4145]; 
    assign out[1870] = layer_0[10557]; 
    assign out[1871] = layer_0[1479]; 
    assign out[1872] = layer_0[3043] ^ layer_0[10594]; 
    assign out[1873] = ~(layer_0[9953] ^ layer_0[5862]); 
    assign out[1874] = ~(layer_0[8189] ^ layer_0[7873]); 
    assign out[1875] = layer_0[2989] & layer_0[9906]; 
    assign out[1876] = layer_0[6952] & ~layer_0[286]; 
    assign out[1877] = layer_0[10249]; 
    assign out[1878] = ~(layer_0[455] ^ layer_0[2292]); 
    assign out[1879] = layer_0[1170] & ~layer_0[3472]; 
    assign out[1880] = ~(layer_0[6133] ^ layer_0[3809]); 
    assign out[1881] = layer_0[1562]; 
    assign out[1882] = layer_0[3513] ^ layer_0[8211]; 
    assign out[1883] = ~(layer_0[564] ^ layer_0[6962]); 
    assign out[1884] = ~(layer_0[2936] ^ layer_0[1107]); 
    assign out[1885] = ~(layer_0[1225] & layer_0[11190]); 
    assign out[1886] = layer_0[6518] & layer_0[10599]; 
    assign out[1887] = layer_0[5383] ^ layer_0[5964]; 
    assign out[1888] = ~layer_0[6965]; 
    assign out[1889] = ~(layer_0[9602] ^ layer_0[2943]); 
    assign out[1890] = layer_0[6320] & layer_0[3822]; 
    assign out[1891] = ~layer_0[3879] | (layer_0[2402] & layer_0[3879]); 
    assign out[1892] = ~(layer_0[5758] ^ layer_0[1278]); 
    assign out[1893] = layer_0[2884] | layer_0[2001]; 
    assign out[1894] = layer_0[1977] ^ layer_0[2501]; 
    assign out[1895] = layer_0[1809] & layer_0[10205]; 
    assign out[1896] = layer_0[10375]; 
    assign out[1897] = ~layer_0[4879]; 
    assign out[1898] = ~(layer_0[2919] ^ layer_0[4708]); 
    assign out[1899] = ~layer_0[6941]; 
    assign out[1900] = layer_0[3502] & ~layer_0[8623]; 
    assign out[1901] = ~layer_0[129]; 
    assign out[1902] = layer_0[4176] ^ layer_0[3564]; 
    assign out[1903] = ~(layer_0[3145] ^ layer_0[4090]); 
    assign out[1904] = layer_0[7216] & ~layer_0[10430]; 
    assign out[1905] = layer_0[1821] ^ layer_0[7822]; 
    assign out[1906] = layer_0[11584] ^ layer_0[4643]; 
    assign out[1907] = ~(layer_0[1481] ^ layer_0[4184]); 
    assign out[1908] = ~(layer_0[7685] ^ layer_0[5624]); 
    assign out[1909] = layer_0[3883] & layer_0[6508]; 
    assign out[1910] = ~(layer_0[1517] ^ layer_0[3781]); 
    assign out[1911] = layer_0[1231] & ~layer_0[7740]; 
    assign out[1912] = ~(layer_0[5665] | layer_0[6580]); 
    assign out[1913] = layer_0[2472] ^ layer_0[11648]; 
    assign out[1914] = layer_0[8657] ^ layer_0[3860]; 
    assign out[1915] = ~(layer_0[4546] ^ layer_0[4924]); 
    assign out[1916] = ~layer_0[9477] | (layer_0[9477] & layer_0[11792]); 
    assign out[1917] = layer_0[1686] & ~layer_0[4974]; 
    assign out[1918] = layer_0[3355] ^ layer_0[10121]; 
    assign out[1919] = ~(layer_0[7472] & layer_0[5744]); 
    assign out[1920] = ~(layer_0[2188] ^ layer_0[4083]); 
    assign out[1921] = layer_0[7339] ^ layer_0[1219]; 
    assign out[1922] = layer_0[1690] ^ layer_0[11797]; 
    assign out[1923] = layer_0[2590] & ~layer_0[2375]; 
    assign out[1924] = layer_0[3400]; 
    assign out[1925] = ~(layer_0[11296] ^ layer_0[9261]); 
    assign out[1926] = layer_0[7241] ^ layer_0[160]; 
    assign out[1927] = layer_0[2846] | layer_0[10896]; 
    assign out[1928] = layer_0[6716] ^ layer_0[7660]; 
    assign out[1929] = ~(layer_0[6857] | layer_0[4572]); 
    assign out[1930] = ~(layer_0[7765] ^ layer_0[2857]); 
    assign out[1931] = layer_0[2497] ^ layer_0[7978]; 
    assign out[1932] = ~(layer_0[8972] & layer_0[7906]); 
    assign out[1933] = ~(layer_0[6346] ^ layer_0[6056]); 
    assign out[1934] = layer_0[9641]; 
    assign out[1935] = ~(layer_0[585] ^ layer_0[683]); 
    assign out[1936] = layer_0[4663] ^ layer_0[5809]; 
    assign out[1937] = layer_0[6760] ^ layer_0[3535]; 
    assign out[1938] = layer_0[6004] ^ layer_0[8151]; 
    assign out[1939] = ~(layer_0[9792] & layer_0[6468]); 
    assign out[1940] = layer_0[6551] & ~layer_0[8917]; 
    assign out[1941] = ~(layer_0[8419] ^ layer_0[7922]); 
    assign out[1942] = ~(layer_0[388] | layer_0[2290]); 
    assign out[1943] = layer_0[3259] & ~layer_0[10173]; 
    assign out[1944] = layer_0[10774] ^ layer_0[7677]; 
    assign out[1945] = layer_0[8610]; 
    assign out[1946] = layer_0[9860] ^ layer_0[212]; 
    assign out[1947] = ~(layer_0[6525] & layer_0[4935]); 
    assign out[1948] = ~(layer_0[3509] ^ layer_0[9929]); 
    assign out[1949] = layer_0[11087] ^ layer_0[7730]; 
    assign out[1950] = layer_0[4120]; 
    assign out[1951] = layer_0[9523] ^ layer_0[1283]; 
    assign out[1952] = ~(layer_0[801] ^ layer_0[3706]); 
    assign out[1953] = layer_0[10038] & ~layer_0[5220]; 
    assign out[1954] = layer_0[9533]; 
    assign out[1955] = layer_0[5528] ^ layer_0[2848]; 
    assign out[1956] = ~layer_0[1892]; 
    assign out[1957] = layer_0[438] & ~layer_0[11751]; 
    assign out[1958] = ~(layer_0[3510] ^ layer_0[7228]); 
    assign out[1959] = ~layer_0[11889]; 
    assign out[1960] = ~(layer_0[11924] ^ layer_0[8730]); 
    assign out[1961] = ~layer_0[1578]; 
    assign out[1962] = layer_0[0] ^ layer_0[5839]; 
    assign out[1963] = ~(layer_0[1728] ^ layer_0[10454]); 
    assign out[1964] = ~(layer_0[294] ^ layer_0[8694]); 
    assign out[1965] = layer_0[8825] ^ layer_0[2607]; 
    assign out[1966] = layer_0[4918] ^ layer_0[3392]; 
    assign out[1967] = ~layer_0[10327]; 
    assign out[1968] = layer_0[6384] ^ layer_0[2306]; 
    assign out[1969] = layer_0[8556] | layer_0[2055]; 
    assign out[1970] = ~layer_0[6220]; 
    assign out[1971] = ~layer_0[1652]; 
    assign out[1972] = layer_0[6216] ^ layer_0[6442]; 
    assign out[1973] = ~layer_0[5906] | (layer_0[4152] & layer_0[5906]); 
    assign out[1974] = ~(layer_0[5141] | layer_0[7963]); 
    assign out[1975] = layer_0[1529] & layer_0[10908]; 
    assign out[1976] = ~layer_0[3011]; 
    assign out[1977] = layer_0[1512]; 
    assign out[1978] = ~(layer_0[6988] ^ layer_0[10799]); 
    assign out[1979] = layer_0[8492] ^ layer_0[8740]; 
    assign out[1980] = layer_0[4071] & layer_0[9252]; 
    assign out[1981] = ~(layer_0[131] ^ layer_0[4011]); 
    assign out[1982] = layer_0[10175] ^ layer_0[7137]; 
    assign out[1983] = layer_0[11781] & ~layer_0[9268]; 
    assign out[1984] = layer_0[444]; 
    assign out[1985] = ~layer_0[2636]; 
    assign out[1986] = layer_0[7093] ^ layer_0[810]; 
    assign out[1987] = ~(layer_0[2737] ^ layer_0[4695]); 
    assign out[1988] = layer_0[1817] ^ layer_0[8073]; 
    assign out[1989] = layer_0[6473] | layer_0[4083]; 
    assign out[1990] = layer_0[11446] & layer_0[6047]; 
    assign out[1991] = layer_0[2235] ^ layer_0[5897]; 
    assign out[1992] = layer_0[1651] & ~layer_0[2514]; 
    assign out[1993] = ~(layer_0[8] ^ layer_0[1418]); 
    assign out[1994] = ~(layer_0[11125] ^ layer_0[3225]); 
    assign out[1995] = ~(layer_0[2635] ^ layer_0[6180]); 
    assign out[1996] = layer_0[11785] ^ layer_0[3350]; 
    assign out[1997] = layer_0[10247] ^ layer_0[8955]; 
    assign out[1998] = ~(layer_0[10752] ^ layer_0[826]); 
    assign out[1999] = layer_0[11039] ^ layer_0[1089]; 
    assign out[2000] = layer_0[7323] & ~layer_0[4934]; 
    assign out[2001] = layer_0[2926] ^ layer_0[1148]; 
    assign out[2002] = ~layer_0[6467]; 
    assign out[2003] = layer_0[11861]; 
    assign out[2004] = layer_0[8301] ^ layer_0[9375]; 
    assign out[2005] = layer_0[11795] ^ layer_0[11366]; 
    assign out[2006] = layer_0[10849]; 
    assign out[2007] = layer_0[6592] ^ layer_0[9558]; 
    assign out[2008] = layer_0[4110] ^ layer_0[2249]; 
    assign out[2009] = ~(layer_0[2066] ^ layer_0[1132]); 
    assign out[2010] = ~(layer_0[2650] ^ layer_0[69]); 
    assign out[2011] = layer_0[7760] ^ layer_0[11375]; 
    assign out[2012] = ~(layer_0[6521] ^ layer_0[9630]); 
    assign out[2013] = ~layer_0[6767]; 
    assign out[2014] = ~layer_0[4030]; 
    assign out[2015] = layer_0[8321] ^ layer_0[5813]; 
    assign out[2016] = layer_0[8508] & ~layer_0[6372]; 
    assign out[2017] = ~(layer_0[7282] ^ layer_0[5316]); 
    assign out[2018] = ~layer_0[9341]; 
    assign out[2019] = ~(layer_0[11981] ^ layer_0[8685]); 
    assign out[2020] = ~(layer_0[2240] ^ layer_0[6412]); 
    assign out[2021] = ~(layer_0[10411] ^ layer_0[4837]); 
    assign out[2022] = layer_0[1737] ^ layer_0[196]; 
    assign out[2023] = layer_0[8286] ^ layer_0[9993]; 
    assign out[2024] = ~(layer_0[7697] ^ layer_0[9601]); 
    assign out[2025] = layer_0[8052] & layer_0[7901]; 
    assign out[2026] = ~(layer_0[10792] | layer_0[4189]); 
    assign out[2027] = ~(layer_0[1221] ^ layer_0[1249]); 
    assign out[2028] = layer_0[4668] & ~layer_0[3483]; 
    assign out[2029] = layer_0[7916] ^ layer_0[6944]; 
    assign out[2030] = layer_0[864] & layer_0[5457]; 
    assign out[2031] = ~(layer_0[4594] ^ layer_0[1932]); 
    assign out[2032] = layer_0[2565] ^ layer_0[11333]; 
    assign out[2033] = layer_0[10817] ^ layer_0[5409]; 
    assign out[2034] = layer_0[560] ^ layer_0[4883]; 
    assign out[2035] = ~(layer_0[4039] ^ layer_0[6833]); 
    assign out[2036] = ~(layer_0[7896] | layer_0[1925]); 
    assign out[2037] = layer_0[5378] ^ layer_0[4514]; 
    assign out[2038] = layer_0[11498] ^ layer_0[9651]; 
    assign out[2039] = ~(layer_0[2390] ^ layer_0[9367]); 
    assign out[2040] = layer_0[8843] & ~layer_0[5515]; 
    assign out[2041] = layer_0[11800] & layer_0[3081]; 
    assign out[2042] = ~(layer_0[11278] ^ layer_0[3842]); 
    assign out[2043] = ~layer_0[314] | (layer_0[5543] & layer_0[314]); 
    assign out[2044] = ~(layer_0[10893] ^ layer_0[6245]); 
    assign out[2045] = ~(layer_0[8629] | layer_0[10233]); 
    assign out[2046] = ~(layer_0[11375] ^ layer_0[3622]); 
    assign out[2047] = ~(layer_0[10068] ^ layer_0[9936]); 
    assign out[2048] = ~layer_0[3786]; 
    assign out[2049] = layer_0[1054]; 
    assign out[2050] = layer_0[4652]; 
    assign out[2051] = ~(layer_0[9833] | layer_0[4010]); 
    assign out[2052] = layer_0[10465] & ~layer_0[5787]; 
    assign out[2053] = layer_0[777] & ~layer_0[57]; 
    assign out[2054] = layer_0[3534] ^ layer_0[4105]; 
    assign out[2055] = ~(layer_0[11825] | layer_0[11439]); 
    assign out[2056] = ~(layer_0[6034] ^ layer_0[4034]); 
    assign out[2057] = layer_0[10312] & ~layer_0[1388]; 
    assign out[2058] = ~(layer_0[1068] | layer_0[174]); 
    assign out[2059] = layer_0[4787] & ~layer_0[1954]; 
    assign out[2060] = layer_0[3560] & ~layer_0[4081]; 
    assign out[2061] = ~(layer_0[11663] ^ layer_0[3948]); 
    assign out[2062] = layer_0[9553] ^ layer_0[1536]; 
    assign out[2063] = layer_0[11880] ^ layer_0[6112]; 
    assign out[2064] = layer_0[6970] ^ layer_0[2839]; 
    assign out[2065] = ~(layer_0[5719] ^ layer_0[7656]); 
    assign out[2066] = layer_0[5894] & layer_0[10275]; 
    assign out[2067] = layer_0[6861] & ~layer_0[11491]; 
    assign out[2068] = layer_0[4866]; 
    assign out[2069] = layer_0[6664]; 
    assign out[2070] = layer_0[4024] & layer_0[2754]; 
    assign out[2071] = ~(layer_0[2217] ^ layer_0[8591]); 
    assign out[2072] = layer_0[335] ^ layer_0[10537]; 
    assign out[2073] = layer_0[1937] ^ layer_0[11717]; 
    assign out[2074] = layer_0[6100] & layer_0[4185]; 
    assign out[2075] = ~layer_0[5575] | (layer_0[10429] & layer_0[5575]); 
    assign out[2076] = layer_0[776] ^ layer_0[232]; 
    assign out[2077] = layer_0[9866] & ~layer_0[6179]; 
    assign out[2078] = ~(layer_0[8470] | layer_0[6003]); 
    assign out[2079] = layer_0[398] & layer_0[5115]; 
    assign out[2080] = ~(layer_0[6915] & layer_0[8997]); 
    assign out[2081] = layer_0[9798] ^ layer_0[10589]; 
    assign out[2082] = layer_0[10528] & ~layer_0[2496]; 
    assign out[2083] = layer_0[5808] & layer_0[8193]; 
    assign out[2084] = ~(layer_0[1560] ^ layer_0[3837]); 
    assign out[2085] = layer_0[5577] | layer_0[7588]; 
    assign out[2086] = layer_0[10024]; 
    assign out[2087] = ~layer_0[7352]; 
    assign out[2088] = ~(layer_0[10489] ^ layer_0[1682]); 
    assign out[2089] = ~(layer_0[1349] ^ layer_0[1428]); 
    assign out[2090] = layer_0[717] & ~layer_0[3311]; 
    assign out[2091] = layer_0[10276] ^ layer_0[7037]; 
    assign out[2092] = ~layer_0[9799]; 
    assign out[2093] = ~layer_0[8219]; 
    assign out[2094] = ~(layer_0[369] ^ layer_0[7867]); 
    assign out[2095] = ~(layer_0[1304] ^ layer_0[4043]); 
    assign out[2096] = ~(layer_0[3095] ^ layer_0[4745]); 
    assign out[2097] = layer_0[10220] ^ layer_0[6343]; 
    assign out[2098] = ~(layer_0[4658] ^ layer_0[11147]); 
    assign out[2099] = ~(layer_0[8352] ^ layer_0[789]); 
    assign out[2100] = layer_0[2286]; 
    assign out[2101] = layer_0[2138]; 
    assign out[2102] = ~layer_0[6832]; 
    assign out[2103] = ~layer_0[3324]; 
    assign out[2104] = ~(layer_0[11195] ^ layer_0[679]); 
    assign out[2105] = layer_0[4068] & ~layer_0[3420]; 
    assign out[2106] = layer_0[6030] & layer_0[4858]; 
    assign out[2107] = layer_0[4950] ^ layer_0[11233]; 
    assign out[2108] = layer_0[6058] & layer_0[4826]; 
    assign out[2109] = ~(layer_0[925] ^ layer_0[4865]); 
    assign out[2110] = ~(layer_0[2045] ^ layer_0[549]); 
    assign out[2111] = layer_0[7271] & ~layer_0[8178]; 
    assign out[2112] = layer_0[558]; 
    assign out[2113] = layer_0[9443] & layer_0[7169]; 
    assign out[2114] = ~(layer_0[9207] ^ layer_0[3485]); 
    assign out[2115] = layer_0[10363] ^ layer_0[7634]; 
    assign out[2116] = layer_0[2676] ^ layer_0[698]; 
    assign out[2117] = ~(layer_0[9207] ^ layer_0[870]); 
    assign out[2118] = ~layer_0[5486]; 
    assign out[2119] = ~(layer_0[2621] | layer_0[10058]); 
    assign out[2120] = layer_0[3359] ^ layer_0[7725]; 
    assign out[2121] = layer_0[5477] & ~layer_0[10058]; 
    assign out[2122] = layer_0[3698] & ~layer_0[9811]; 
    assign out[2123] = ~layer_0[4912]; 
    assign out[2124] = ~(layer_0[1556] ^ layer_0[4143]); 
    assign out[2125] = ~(layer_0[2784] | layer_0[5176]); 
    assign out[2126] = layer_0[2377] & ~layer_0[1243]; 
    assign out[2127] = layer_0[5282]; 
    assign out[2128] = layer_0[7363] ^ layer_0[5388]; 
    assign out[2129] = ~layer_0[3728]; 
    assign out[2130] = layer_0[1979]; 
    assign out[2131] = ~(layer_0[10200] ^ layer_0[6110]); 
    assign out[2132] = layer_0[7698] ^ layer_0[6636]; 
    assign out[2133] = ~(layer_0[3403] ^ layer_0[171]); 
    assign out[2134] = layer_0[8792] ^ layer_0[688]; 
    assign out[2135] = ~(layer_0[9029] ^ layer_0[3533]); 
    assign out[2136] = layer_0[5424] | layer_0[4901]; 
    assign out[2137] = layer_0[6093] ^ layer_0[9657]; 
    assign out[2138] = layer_0[7827] ^ layer_0[8389]; 
    assign out[2139] = ~(layer_0[10853] ^ layer_0[7328]); 
    assign out[2140] = layer_0[7246]; 
    assign out[2141] = layer_0[10311] ^ layer_0[8976]; 
    assign out[2142] = ~(layer_0[9633] | layer_0[1845]); 
    assign out[2143] = ~(layer_0[4154] ^ layer_0[6887]); 
    assign out[2144] = ~(layer_0[10777] ^ layer_0[8975]); 
    assign out[2145] = ~(layer_0[1261] ^ layer_0[8450]); 
    assign out[2146] = ~(layer_0[1368] ^ layer_0[3953]); 
    assign out[2147] = ~layer_0[10418] | (layer_0[4279] & layer_0[10418]); 
    assign out[2148] = layer_0[674]; 
    assign out[2149] = ~(layer_0[4519] ^ layer_0[7716]); 
    assign out[2150] = ~(layer_0[7222] ^ layer_0[2765]); 
    assign out[2151] = ~layer_0[9234] | (layer_0[5272] & layer_0[9234]); 
    assign out[2152] = ~layer_0[11873]; 
    assign out[2153] = layer_0[2639] ^ layer_0[147]; 
    assign out[2154] = layer_0[5313] | layer_0[9935]; 
    assign out[2155] = layer_0[1657]; 
    assign out[2156] = ~(layer_0[3079] ^ layer_0[9785]); 
    assign out[2157] = layer_0[7922] | layer_0[11021]; 
    assign out[2158] = layer_0[6764] ^ layer_0[7783]; 
    assign out[2159] = ~(layer_0[9249] ^ layer_0[8444]); 
    assign out[2160] = layer_0[11882] | layer_0[4891]; 
    assign out[2161] = ~(layer_0[3950] ^ layer_0[6308]); 
    assign out[2162] = layer_0[11696] ^ layer_0[7598]; 
    assign out[2163] = layer_0[4366] & layer_0[11]; 
    assign out[2164] = ~(layer_0[1961] ^ layer_0[3918]); 
    assign out[2165] = layer_0[4065] ^ layer_0[3906]; 
    assign out[2166] = ~(layer_0[11076] ^ layer_0[9400]); 
    assign out[2167] = layer_0[3257] & ~layer_0[5501]; 
    assign out[2168] = ~layer_0[8261]; 
    assign out[2169] = layer_0[7891] ^ layer_0[4601]; 
    assign out[2170] = ~(layer_0[2866] ^ layer_0[1955]); 
    assign out[2171] = layer_0[41] & ~layer_0[2195]; 
    assign out[2172] = layer_0[2488] ^ layer_0[2804]; 
    assign out[2173] = ~layer_0[6487]; 
    assign out[2174] = ~(layer_0[6930] ^ layer_0[6295]); 
    assign out[2175] = ~(layer_0[9049] ^ layer_0[9948]); 
    assign out[2176] = ~(layer_0[11996] ^ layer_0[11533]); 
    assign out[2177] = layer_0[1384]; 
    assign out[2178] = ~layer_0[35]; 
    assign out[2179] = ~(layer_0[10732] ^ layer_0[353]); 
    assign out[2180] = ~(layer_0[10195] ^ layer_0[3210]); 
    assign out[2181] = ~(layer_0[852] ^ layer_0[2526]); 
    assign out[2182] = ~(layer_0[117] ^ layer_0[4856]); 
    assign out[2183] = layer_0[9818] ^ layer_0[877]; 
    assign out[2184] = layer_0[10336] & layer_0[111]; 
    assign out[2185] = ~(layer_0[2399] ^ layer_0[8050]); 
    assign out[2186] = ~(layer_0[4794] & layer_0[8423]); 
    assign out[2187] = ~(layer_0[3891] ^ layer_0[3479]); 
    assign out[2188] = layer_0[5919] ^ layer_0[3809]; 
    assign out[2189] = ~layer_0[1145] | (layer_0[3387] & layer_0[1145]); 
    assign out[2190] = layer_0[4873] & layer_0[4588]; 
    assign out[2191] = ~(layer_0[4331] & layer_0[3911]); 
    assign out[2192] = layer_0[3261]; 
    assign out[2193] = layer_0[1869] ^ layer_0[2922]; 
    assign out[2194] = ~(layer_0[3363] ^ layer_0[3999]); 
    assign out[2195] = layer_0[2629] ^ layer_0[3763]; 
    assign out[2196] = ~(layer_0[10143] | layer_0[9047]); 
    assign out[2197] = ~(layer_0[5268] ^ layer_0[8750]); 
    assign out[2198] = layer_0[4923] ^ layer_0[1940]; 
    assign out[2199] = layer_0[10728] ^ layer_0[6423]; 
    assign out[2200] = ~(layer_0[11153] ^ layer_0[3435]); 
    assign out[2201] = layer_0[6166] ^ layer_0[2002]; 
    assign out[2202] = ~(layer_0[3743] ^ layer_0[714]); 
    assign out[2203] = layer_0[6730] ^ layer_0[10529]; 
    assign out[2204] = ~(layer_0[6593] ^ layer_0[3767]); 
    assign out[2205] = ~layer_0[3341] | (layer_0[3341] & layer_0[3443]); 
    assign out[2206] = ~(layer_0[4841] ^ layer_0[4916]); 
    assign out[2207] = ~(layer_0[10413] ^ layer_0[11062]); 
    assign out[2208] = ~layer_0[5890] | (layer_0[5510] & layer_0[5890]); 
    assign out[2209] = layer_0[8006] ^ layer_0[8795]; 
    assign out[2210] = ~(layer_0[6119] | layer_0[11341]); 
    assign out[2211] = layer_0[8516] ^ layer_0[6945]; 
    assign out[2212] = layer_0[5873] ^ layer_0[170]; 
    assign out[2213] = layer_0[3926] | layer_0[4310]; 
    assign out[2214] = layer_0[2232] ^ layer_0[5010]; 
    assign out[2215] = layer_0[10562] ^ layer_0[4733]; 
    assign out[2216] = ~(layer_0[10435] | layer_0[4502]); 
    assign out[2217] = layer_0[9406] | layer_0[475]; 
    assign out[2218] = layer_0[8583] & ~layer_0[6788]; 
    assign out[2219] = layer_0[9067] ^ layer_0[8592]; 
    assign out[2220] = layer_0[6117]; 
    assign out[2221] = layer_0[7223] ^ layer_0[7610]; 
    assign out[2222] = layer_0[6330] ^ layer_0[2790]; 
    assign out[2223] = ~(layer_0[10788] ^ layer_0[957]); 
    assign out[2224] = ~(layer_0[4032] ^ layer_0[7382]); 
    assign out[2225] = ~(layer_0[2927] ^ layer_0[8669]); 
    assign out[2226] = layer_0[10843]; 
    assign out[2227] = layer_0[726] ^ layer_0[9095]; 
    assign out[2228] = layer_0[4289] ^ layer_0[2128]; 
    assign out[2229] = layer_0[10926] ^ layer_0[5613]; 
    assign out[2230] = ~(layer_0[5104] ^ layer_0[10671]); 
    assign out[2231] = layer_0[4427] ^ layer_0[10172]; 
    assign out[2232] = layer_0[5249] ^ layer_0[5869]; 
    assign out[2233] = ~layer_0[1919] | (layer_0[1919] & layer_0[11951]); 
    assign out[2234] = layer_0[2703]; 
    assign out[2235] = layer_0[5926] ^ layer_0[8760]; 
    assign out[2236] = ~layer_0[8182] | (layer_0[8182] & layer_0[1705]); 
    assign out[2237] = layer_0[2709] ^ layer_0[7301]; 
    assign out[2238] = layer_0[9409] ^ layer_0[10667]; 
    assign out[2239] = layer_0[3808] | layer_0[8511]; 
    assign out[2240] = layer_0[3138] ^ layer_0[6946]; 
    assign out[2241] = layer_0[4807] ^ layer_0[2575]; 
    assign out[2242] = layer_0[1311] ^ layer_0[4899]; 
    assign out[2243] = layer_0[8006] & ~layer_0[7585]; 
    assign out[2244] = layer_0[5696] & layer_0[7671]; 
    assign out[2245] = ~(layer_0[5279] ^ layer_0[126]); 
    assign out[2246] = ~layer_0[10988]; 
    assign out[2247] = ~layer_0[8768]; 
    assign out[2248] = ~(layer_0[3495] & layer_0[843]); 
    assign out[2249] = ~(layer_0[10097] ^ layer_0[11748]); 
    assign out[2250] = ~(layer_0[10754] ^ layer_0[8745]); 
    assign out[2251] = layer_0[7681] & layer_0[8518]; 
    assign out[2252] = ~(layer_0[5632] ^ layer_0[4651]); 
    assign out[2253] = layer_0[248] & ~layer_0[9191]; 
    assign out[2254] = layer_0[3286] & layer_0[7704]; 
    assign out[2255] = layer_0[555] & layer_0[1474]; 
    assign out[2256] = layer_0[2274] & ~layer_0[5300]; 
    assign out[2257] = ~(layer_0[10576] | layer_0[11225]); 
    assign out[2258] = ~(layer_0[1770] ^ layer_0[11647]); 
    assign out[2259] = ~(layer_0[11761] | layer_0[1884]); 
    assign out[2260] = ~layer_0[1799]; 
    assign out[2261] = ~layer_0[923] | (layer_0[5532] & layer_0[923]); 
    assign out[2262] = layer_0[9620] | layer_0[7941]; 
    assign out[2263] = layer_0[11983] & ~layer_0[11741]; 
    assign out[2264] = layer_0[3952] ^ layer_0[8944]; 
    assign out[2265] = ~(layer_0[3273] | layer_0[6961]); 
    assign out[2266] = layer_0[5078]; 
    assign out[2267] = ~layer_0[4407]; 
    assign out[2268] = layer_0[6548]; 
    assign out[2269] = layer_0[5746] ^ layer_0[2270]; 
    assign out[2270] = layer_0[2774] & ~layer_0[11221]; 
    assign out[2271] = layer_0[1003] ^ layer_0[11336]; 
    assign out[2272] = layer_0[10737]; 
    assign out[2273] = layer_0[394] ^ layer_0[3012]; 
    assign out[2274] = layer_0[3796] & ~layer_0[10643]; 
    assign out[2275] = layer_0[1047] ^ layer_0[10804]; 
    assign out[2276] = ~layer_0[5225]; 
    assign out[2277] = ~layer_0[10504]; 
    assign out[2278] = ~(layer_0[6264] ^ layer_0[2484]); 
    assign out[2279] = ~layer_0[8940]; 
    assign out[2280] = layer_0[8527] & ~layer_0[10468]; 
    assign out[2281] = ~(layer_0[11934] | layer_0[3222]); 
    assign out[2282] = ~(layer_0[11949] ^ layer_0[10918]); 
    assign out[2283] = ~layer_0[5552] | (layer_0[9914] & layer_0[5552]); 
    assign out[2284] = layer_0[4993] ^ layer_0[2230]; 
    assign out[2285] = ~(layer_0[8371] & layer_0[205]); 
    assign out[2286] = layer_0[7445]; 
    assign out[2287] = ~(layer_0[8175] ^ layer_0[3040]); 
    assign out[2288] = layer_0[10821] & ~layer_0[9454]; 
    assign out[2289] = ~(layer_0[5126] | layer_0[6910]); 
    assign out[2290] = layer_0[7823] ^ layer_0[8132]; 
    assign out[2291] = layer_0[1096] & ~layer_0[1283]; 
    assign out[2292] = ~(layer_0[3425] & layer_0[7999]); 
    assign out[2293] = layer_0[10507] & ~layer_0[10378]; 
    assign out[2294] = ~(layer_0[4959] & layer_0[11594]); 
    assign out[2295] = layer_0[11983] & ~layer_0[3605]; 
    assign out[2296] = layer_0[409] ^ layer_0[7869]; 
    assign out[2297] = layer_0[6064] | layer_0[3366]; 
    assign out[2298] = layer_0[344]; 
    assign out[2299] = layer_0[2813] ^ layer_0[4876]; 
    assign out[2300] = ~(layer_0[4876] ^ layer_0[1577]); 
    assign out[2301] = layer_0[10908]; 
    assign out[2302] = ~layer_0[9746]; 
    assign out[2303] = ~(layer_0[4046] ^ layer_0[10920]); 
    assign out[2304] = ~layer_0[11865]; 
    assign out[2305] = ~(layer_0[1936] ^ layer_0[10033]); 
    assign out[2306] = layer_0[4942] & ~layer_0[11836]; 
    assign out[2307] = ~(layer_0[11691] | layer_0[2771]); 
    assign out[2308] = ~(layer_0[2555] ^ layer_0[7820]); 
    assign out[2309] = layer_0[4496] ^ layer_0[11947]; 
    assign out[2310] = layer_0[9366] ^ layer_0[4877]; 
    assign out[2311] = layer_0[11095] | layer_0[8709]; 
    assign out[2312] = ~layer_0[4177]; 
    assign out[2313] = ~(layer_0[10402] ^ layer_0[5715]); 
    assign out[2314] = layer_0[4612] ^ layer_0[7132]; 
    assign out[2315] = layer_0[11457] & layer_0[11284]; 
    assign out[2316] = layer_0[9471] & ~layer_0[1183]; 
    assign out[2317] = layer_0[10317]; 
    assign out[2318] = ~(layer_0[7118] ^ layer_0[6377]); 
    assign out[2319] = ~(layer_0[7142] ^ layer_0[2545]); 
    assign out[2320] = ~(layer_0[3115] ^ layer_0[1041]); 
    assign out[2321] = layer_0[8854] ^ layer_0[10370]; 
    assign out[2322] = layer_0[9337]; 
    assign out[2323] = layer_0[8995] ^ layer_0[10064]; 
    assign out[2324] = layer_0[1528] ^ layer_0[3369]; 
    assign out[2325] = ~layer_0[1189]; 
    assign out[2326] = ~layer_0[11307] | (layer_0[8312] & layer_0[11307]); 
    assign out[2327] = ~(layer_0[2601] ^ layer_0[8923]); 
    assign out[2328] = ~(layer_0[3740] ^ layer_0[2160]); 
    assign out[2329] = layer_0[9346] ^ layer_0[307]; 
    assign out[2330] = ~(layer_0[8325] ^ layer_0[20]); 
    assign out[2331] = ~layer_0[7011] | (layer_0[2147] & layer_0[7011]); 
    assign out[2332] = ~(layer_0[509] | layer_0[3693]); 
    assign out[2333] = layer_0[2219]; 
    assign out[2334] = ~(layer_0[3090] ^ layer_0[5900]); 
    assign out[2335] = layer_0[6464] ^ layer_0[893]; 
    assign out[2336] = layer_0[10692] & layer_0[10003]; 
    assign out[2337] = layer_0[3072]; 
    assign out[2338] = ~layer_0[4744]; 
    assign out[2339] = layer_0[2662] & layer_0[710]; 
    assign out[2340] = layer_0[7247] ^ layer_0[4106]; 
    assign out[2341] = ~layer_0[8787]; 
    assign out[2342] = ~layer_0[1408]; 
    assign out[2343] = ~(layer_0[987] ^ layer_0[7406]); 
    assign out[2344] = ~(layer_0[11993] | layer_0[1255]); 
    assign out[2345] = ~(layer_0[4872] ^ layer_0[1775]); 
    assign out[2346] = layer_0[10882] | layer_0[11334]; 
    assign out[2347] = ~(layer_0[4130] ^ layer_0[9091]); 
    assign out[2348] = layer_0[2208] ^ layer_0[11837]; 
    assign out[2349] = layer_0[9563]; 
    assign out[2350] = layer_0[740] ^ layer_0[4429]; 
    assign out[2351] = layer_0[8252] & ~layer_0[603]; 
    assign out[2352] = ~(layer_0[10828] ^ layer_0[9578]); 
    assign out[2353] = layer_0[6747] ^ layer_0[3473]; 
    assign out[2354] = layer_0[1045] ^ layer_0[6088]; 
    assign out[2355] = ~layer_0[4983] | (layer_0[4983] & layer_0[2474]); 
    assign out[2356] = layer_0[9407] & ~layer_0[1376]; 
    assign out[2357] = layer_0[1893] ^ layer_0[2971]; 
    assign out[2358] = layer_0[835]; 
    assign out[2359] = ~(layer_0[6140] ^ layer_0[7059]); 
    assign out[2360] = layer_0[7356] ^ layer_0[2061]; 
    assign out[2361] = ~(layer_0[7192] ^ layer_0[3886]); 
    assign out[2362] = ~layer_0[4502]; 
    assign out[2363] = ~layer_0[9895] | (layer_0[9895] & layer_0[7610]); 
    assign out[2364] = layer_0[2895] & ~layer_0[752]; 
    assign out[2365] = layer_0[9764] & layer_0[10599]; 
    assign out[2366] = layer_0[1752]; 
    assign out[2367] = ~(layer_0[1418] ^ layer_0[543]); 
    assign out[2368] = layer_0[9910] ^ layer_0[7976]; 
    assign out[2369] = layer_0[6501]; 
    assign out[2370] = ~(layer_0[5399] ^ layer_0[4220]); 
    assign out[2371] = ~(layer_0[4016] ^ layer_0[8065]); 
    assign out[2372] = ~(layer_0[3348] ^ layer_0[7324]); 
    assign out[2373] = layer_0[10302]; 
    assign out[2374] = ~layer_0[8783]; 
    assign out[2375] = layer_0[1746]; 
    assign out[2376] = ~(layer_0[2336] | layer_0[6303]); 
    assign out[2377] = layer_0[6307] & layer_0[4230]; 
    assign out[2378] = layer_0[1113]; 
    assign out[2379] = layer_0[4820] ^ layer_0[2975]; 
    assign out[2380] = layer_0[1734] ^ layer_0[7943]; 
    assign out[2381] = layer_0[7355] & layer_0[7097]; 
    assign out[2382] = ~(layer_0[8651] ^ layer_0[8452]); 
    assign out[2383] = layer_0[2696] ^ layer_0[10720]; 
    assign out[2384] = layer_0[4277]; 
    assign out[2385] = layer_0[83]; 
    assign out[2386] = ~(layer_0[7145] & layer_0[11247]); 
    assign out[2387] = layer_0[5410]; 
    assign out[2388] = ~(layer_0[10134] ^ layer_0[11394]); 
    assign out[2389] = layer_0[10740] ^ layer_0[6890]; 
    assign out[2390] = layer_0[2930] ^ layer_0[8263]; 
    assign out[2391] = layer_0[11428] ^ layer_0[11087]; 
    assign out[2392] = ~(layer_0[11014] ^ layer_0[8980]); 
    assign out[2393] = ~(layer_0[10567] ^ layer_0[2724]); 
    assign out[2394] = layer_0[8353] & layer_0[1890]; 
    assign out[2395] = layer_0[3653] ^ layer_0[1056]; 
    assign out[2396] = ~(layer_0[621] ^ layer_0[6892]); 
    assign out[2397] = layer_0[4969]; 
    assign out[2398] = ~(layer_0[5616] | layer_0[3907]); 
    assign out[2399] = ~(layer_0[1081] ^ layer_0[451]); 
    assign out[2400] = layer_0[10974] ^ layer_0[5611]; 
    assign out[2401] = ~(layer_0[10360] ^ layer_0[8550]); 
    assign out[2402] = layer_0[2301]; 
    assign out[2403] = layer_0[6859] & ~layer_0[4141]; 
    assign out[2404] = ~(layer_0[7773] ^ layer_0[11373]); 
    assign out[2405] = layer_0[5381] ^ layer_0[5704]; 
    assign out[2406] = ~(layer_0[2979] ^ layer_0[2862]); 
    assign out[2407] = layer_0[6113] | layer_0[9134]; 
    assign out[2408] = layer_0[3062] & ~layer_0[10383]; 
    assign out[2409] = ~layer_0[10544]; 
    assign out[2410] = layer_0[5485] ^ layer_0[8470]; 
    assign out[2411] = ~layer_0[6431]; 
    assign out[2412] = ~(layer_0[4995] ^ layer_0[3426]); 
    assign out[2413] = layer_0[6524]; 
    assign out[2414] = layer_0[10132] & ~layer_0[11869]; 
    assign out[2415] = layer_0[4691] ^ layer_0[1705]; 
    assign out[2416] = ~(layer_0[6364] ^ layer_0[8467]); 
    assign out[2417] = layer_0[3908] & layer_0[463]; 
    assign out[2418] = ~layer_0[3575]; 
    assign out[2419] = ~(layer_0[5432] ^ layer_0[213]); 
    assign out[2420] = layer_0[4793] ^ layer_0[5707]; 
    assign out[2421] = layer_0[7308] ^ layer_0[11040]; 
    assign out[2422] = layer_0[1006] ^ layer_0[6564]; 
    assign out[2423] = ~(layer_0[450] ^ layer_0[1174]); 
    assign out[2424] = ~(layer_0[11312] | layer_0[6523]); 
    assign out[2425] = layer_0[2315] ^ layer_0[1110]; 
    assign out[2426] = ~(layer_0[4766] ^ layer_0[1217]); 
    assign out[2427] = ~(layer_0[2877] ^ layer_0[11679]); 
    assign out[2428] = ~(layer_0[2373] | layer_0[2482]); 
    assign out[2429] = ~(layer_0[7227] | layer_0[9707]); 
    assign out[2430] = layer_0[9600] & ~layer_0[5361]; 
    assign out[2431] = layer_0[3379] ^ layer_0[7510]; 
    assign out[2432] = layer_0[11560] ^ layer_0[3042]; 
    assign out[2433] = layer_0[5042] & ~layer_0[6711]; 
    assign out[2434] = ~(layer_0[7957] ^ layer_0[2661]); 
    assign out[2435] = layer_0[4957] ^ layer_0[1329]; 
    assign out[2436] = layer_0[10406] ^ layer_0[11933]; 
    assign out[2437] = ~layer_0[5957] | (layer_0[5957] & layer_0[9381]); 
    assign out[2438] = ~(layer_0[2981] ^ layer_0[11077]); 
    assign out[2439] = ~layer_0[5989] | (layer_0[8210] & layer_0[5989]); 
    assign out[2440] = layer_0[6869] ^ layer_0[7696]; 
    assign out[2441] = layer_0[8532] | layer_0[894]; 
    assign out[2442] = layer_0[11048] ^ layer_0[1545]; 
    assign out[2443] = ~(layer_0[8106] ^ layer_0[2291]); 
    assign out[2444] = layer_0[6198] ^ layer_0[8152]; 
    assign out[2445] = ~(layer_0[7183] ^ layer_0[625]); 
    assign out[2446] = layer_0[7346] ^ layer_0[11138]; 
    assign out[2447] = ~layer_0[8998] | (layer_0[8998] & layer_0[1475]); 
    assign out[2448] = ~(layer_0[5921] ^ layer_0[5756]); 
    assign out[2449] = layer_0[5572] & ~layer_0[11086]; 
    assign out[2450] = layer_0[6709] ^ layer_0[10069]; 
    assign out[2451] = layer_0[3423] ^ layer_0[5693]; 
    assign out[2452] = layer_0[5891]; 
    assign out[2453] = ~(layer_0[4988] ^ layer_0[6101]); 
    assign out[2454] = layer_0[3684] | layer_0[7369]; 
    assign out[2455] = layer_0[9955] ^ layer_0[6810]; 
    assign out[2456] = ~(layer_0[8534] ^ layer_0[4264]); 
    assign out[2457] = layer_0[2442] ^ layer_0[1164]; 
    assign out[2458] = ~layer_0[4967] | (layer_0[2943] & layer_0[4967]); 
    assign out[2459] = layer_0[7609] & ~layer_0[560]; 
    assign out[2460] = ~(layer_0[180] | layer_0[1156]); 
    assign out[2461] = ~(layer_0[10891] & layer_0[9376]); 
    assign out[2462] = layer_0[10186] ^ layer_0[8775]; 
    assign out[2463] = ~(layer_0[8700] | layer_0[755]); 
    assign out[2464] = layer_0[8310] & ~layer_0[93]; 
    assign out[2465] = ~(layer_0[5747] ^ layer_0[7813]); 
    assign out[2466] = layer_0[2413] ^ layer_0[1486]; 
    assign out[2467] = layer_0[11695]; 
    assign out[2468] = layer_0[7024] & ~layer_0[7990]; 
    assign out[2469] = layer_0[9884] ^ layer_0[7502]; 
    assign out[2470] = ~(layer_0[10256] ^ layer_0[8003]); 
    assign out[2471] = ~layer_0[2694]; 
    assign out[2472] = ~(layer_0[4532] & layer_0[3603]); 
    assign out[2473] = layer_0[1467] & ~layer_0[8593]; 
    assign out[2474] = layer_0[7025] ^ layer_0[487]; 
    assign out[2475] = layer_0[7724] ^ layer_0[11583]; 
    assign out[2476] = layer_0[4271]; 
    assign out[2477] = ~(layer_0[24] | layer_0[7877]); 
    assign out[2478] = ~(layer_0[9711] ^ layer_0[8164]); 
    assign out[2479] = layer_0[9212] & ~layer_0[9743]; 
    assign out[2480] = ~(layer_0[5939] ^ layer_0[5518]); 
    assign out[2481] = ~layer_0[1415]; 
    assign out[2482] = layer_0[3627] | layer_0[1455]; 
    assign out[2483] = layer_0[7767]; 
    assign out[2484] = layer_0[4256] ^ layer_0[5308]; 
    assign out[2485] = ~(layer_0[1997] ^ layer_0[8801]); 
    assign out[2486] = ~(layer_0[10149] | layer_0[8643]); 
    assign out[2487] = layer_0[9065] ^ layer_0[9224]; 
    assign out[2488] = ~(layer_0[558] ^ layer_0[2213]); 
    assign out[2489] = layer_0[6466] & ~layer_0[7587]; 
    assign out[2490] = ~(layer_0[2129] ^ layer_0[8487]); 
    assign out[2491] = layer_0[1394] ^ layer_0[76]; 
    assign out[2492] = layer_0[10184] ^ layer_0[3290]; 
    assign out[2493] = ~(layer_0[11957] ^ layer_0[5496]); 
    assign out[2494] = ~layer_0[3019]; 
    assign out[2495] = ~(layer_0[6642] | layer_0[8337]); 
    assign out[2496] = ~(layer_0[1451] | layer_0[335]); 
    assign out[2497] = layer_0[3219] & ~layer_0[1836]; 
    assign out[2498] = ~(layer_0[9323] ^ layer_0[2350]); 
    assign out[2499] = layer_0[7857] ^ layer_0[4183]; 
    assign out[2500] = ~layer_0[7392] | (layer_0[8435] & layer_0[7392]); 
    assign out[2501] = ~(layer_0[8341] ^ layer_0[461]); 
    assign out[2502] = ~(layer_0[263] ^ layer_0[4791]); 
    assign out[2503] = ~(layer_0[3730] ^ layer_0[4075]); 
    assign out[2504] = layer_0[11545]; 
    assign out[2505] = layer_0[7332] ^ layer_0[5237]; 
    assign out[2506] = ~layer_0[8405]; 
    assign out[2507] = layer_0[5810] | layer_0[8268]; 
    assign out[2508] = ~layer_0[400] | (layer_0[400] & layer_0[3234]); 
    assign out[2509] = ~layer_0[2420] | (layer_0[8963] & layer_0[2420]); 
    assign out[2510] = layer_0[8152]; 
    assign out[2511] = ~(layer_0[1147] ^ layer_0[7513]); 
    assign out[2512] = ~(layer_0[8368] ^ layer_0[10658]); 
    assign out[2513] = ~(layer_0[9831] ^ layer_0[7762]); 
    assign out[2514] = layer_0[1720] ^ layer_0[5707]; 
    assign out[2515] = layer_0[9541] ^ layer_0[2907]; 
    assign out[2516] = layer_0[2822]; 
    assign out[2517] = ~(layer_0[10970] ^ layer_0[8831]); 
    assign out[2518] = layer_0[1372] & ~layer_0[1472]; 
    assign out[2519] = ~layer_0[2649] | (layer_0[9007] & layer_0[2649]); 
    assign out[2520] = layer_0[11025] & ~layer_0[10739]; 
    assign out[2521] = layer_0[7866] ^ layer_0[10932]; 
    assign out[2522] = ~layer_0[3915]; 
    assign out[2523] = layer_0[2214] & ~layer_0[3619]; 
    assign out[2524] = ~(layer_0[7020] ^ layer_0[4933]); 
    assign out[2525] = layer_0[1908] & ~layer_0[10924]; 
    assign out[2526] = layer_0[9089]; 
    assign out[2527] = ~layer_0[1669] | (layer_0[1669] & layer_0[1500]); 
    assign out[2528] = layer_0[8824] & layer_0[5853]; 
    assign out[2529] = layer_0[9241] & layer_0[4176]; 
    assign out[2530] = layer_0[8179] ^ layer_0[2982]; 
    assign out[2531] = ~layer_0[623]; 
    assign out[2532] = ~layer_0[6801] | (layer_0[6801] & layer_0[3249]); 
    assign out[2533] = ~layer_0[10773] | (layer_0[7705] & layer_0[10773]); 
    assign out[2534] = ~(layer_0[9863] ^ layer_0[5672]); 
    assign out[2535] = layer_0[2142] ^ layer_0[4131]; 
    assign out[2536] = layer_0[11278] ^ layer_0[4595]; 
    assign out[2537] = layer_0[10772] ^ layer_0[7937]; 
    assign out[2538] = layer_0[2057]; 
    assign out[2539] = ~(layer_0[5109] ^ layer_0[633]); 
    assign out[2540] = ~(layer_0[9512] ^ layer_0[2949]); 
    assign out[2541] = ~layer_0[8759]; 
    assign out[2542] = ~(layer_0[899] | layer_0[3613]); 
    assign out[2543] = ~(layer_0[1679] ^ layer_0[11361]); 
    assign out[2544] = ~(layer_0[4251] & layer_0[10224]); 
    assign out[2545] = layer_0[10524] ^ layer_0[2260]; 
    assign out[2546] = layer_0[6569] ^ layer_0[9618]; 
    assign out[2547] = ~layer_0[5811]; 
    assign out[2548] = ~(layer_0[3258] ^ layer_0[3424]); 
    assign out[2549] = ~(layer_0[11940] ^ layer_0[8166]); 
    assign out[2550] = layer_0[4420] & ~layer_0[3181]; 
    assign out[2551] = layer_0[772] ^ layer_0[8222]; 
    assign out[2552] = ~(layer_0[211] ^ layer_0[8334]); 
    assign out[2553] = ~(layer_0[6965] ^ layer_0[9359]); 
    assign out[2554] = layer_0[6085] | layer_0[1360]; 
    assign out[2555] = layer_0[2775] ^ layer_0[948]; 
    assign out[2556] = ~layer_0[8810]; 
    assign out[2557] = ~(layer_0[8714] ^ layer_0[2480]); 
    assign out[2558] = layer_0[11242] ^ layer_0[5829]; 
    assign out[2559] = layer_0[6509] | layer_0[460]; 
    assign out[2560] = layer_0[5656]; 
    assign out[2561] = layer_0[3771]; 
    assign out[2562] = ~layer_0[7078]; 
    assign out[2563] = layer_0[7445] & ~layer_0[38]; 
    assign out[2564] = ~(layer_0[6104] ^ layer_0[8727]); 
    assign out[2565] = 1'b0; 
    assign out[2566] = layer_0[2889] ^ layer_0[4055]; 
    assign out[2567] = ~(layer_0[11830] | layer_0[8143]); 
    assign out[2568] = layer_0[7207] ^ layer_0[6351]; 
    assign out[2569] = layer_0[10966] ^ layer_0[5310]; 
    assign out[2570] = ~layer_0[377] | (layer_0[377] & layer_0[1146]); 
    assign out[2571] = layer_0[5814]; 
    assign out[2572] = layer_0[11596] ^ layer_0[8092]; 
    assign out[2573] = layer_0[8983]; 
    assign out[2574] = layer_0[11946] & ~layer_0[4838]; 
    assign out[2575] = layer_0[4136] ^ layer_0[1511]; 
    assign out[2576] = ~(layer_0[9853] ^ layer_0[7121]); 
    assign out[2577] = ~(layer_0[5826] ^ layer_0[10906]); 
    assign out[2578] = layer_0[1485] ^ layer_0[10664]; 
    assign out[2579] = ~layer_0[2209] | (layer_0[10272] & layer_0[2209]); 
    assign out[2580] = layer_0[11652]; 
    assign out[2581] = layer_0[9124]; 
    assign out[2582] = ~(layer_0[9077] ^ layer_0[3881]); 
    assign out[2583] = layer_0[7199]; 
    assign out[2584] = ~layer_0[11290]; 
    assign out[2585] = layer_0[1841]; 
    assign out[2586] = layer_0[9085] & ~layer_0[3929]; 
    assign out[2587] = ~layer_0[6381] | (layer_0[6381] & layer_0[9157]); 
    assign out[2588] = layer_0[3285] ^ layer_0[7693]; 
    assign out[2589] = ~layer_0[694]; 
    assign out[2590] = ~(layer_0[4716] & layer_0[7101]); 
    assign out[2591] = ~(layer_0[1655] ^ layer_0[8743]); 
    assign out[2592] = layer_0[915] | layer_0[7974]; 
    assign out[2593] = layer_0[9291] ^ layer_0[2201]; 
    assign out[2594] = ~(layer_0[7404] ^ layer_0[5952]); 
    assign out[2595] = ~(layer_0[5198] ^ layer_0[11738]); 
    assign out[2596] = layer_0[1442] ^ layer_0[11171]; 
    assign out[2597] = layer_0[9717] & layer_0[3429]; 
    assign out[2598] = layer_0[4622] ^ layer_0[7685]; 
    assign out[2599] = ~(layer_0[9466] ^ layer_0[2014]); 
    assign out[2600] = ~layer_0[1405]; 
    assign out[2601] = layer_0[10170] ^ layer_0[1450]; 
    assign out[2602] = layer_0[10936] | layer_0[5394]; 
    assign out[2603] = layer_0[6543] & ~layer_0[2563]; 
    assign out[2604] = layer_0[5159] ^ layer_0[10409]; 
    assign out[2605] = layer_0[1729] | layer_0[8138]; 
    assign out[2606] = layer_0[7268]; 
    assign out[2607] = ~(layer_0[8013] ^ layer_0[212]); 
    assign out[2608] = ~layer_0[3468]; 
    assign out[2609] = layer_0[11529]; 
    assign out[2610] = layer_0[6399] & ~layer_0[8040]; 
    assign out[2611] = layer_0[8324]; 
    assign out[2612] = ~(layer_0[9342] ^ layer_0[6729]); 
    assign out[2613] = layer_0[9645] ^ layer_0[9281]; 
    assign out[2614] = layer_0[3289] ^ layer_0[10860]; 
    assign out[2615] = ~(layer_0[2551] ^ layer_0[3847]); 
    assign out[2616] = layer_0[8912] ^ layer_0[6211]; 
    assign out[2617] = layer_0[5286] | layer_0[11698]; 
    assign out[2618] = layer_0[9591] & ~layer_0[5990]; 
    assign out[2619] = ~(layer_0[46] ^ layer_0[4864]); 
    assign out[2620] = ~(layer_0[2860] | layer_0[655]); 
    assign out[2621] = layer_0[10928] ^ layer_0[8957]; 
    assign out[2622] = layer_0[2529] & ~layer_0[2746]; 
    assign out[2623] = layer_0[5691] & ~layer_0[8768]; 
    assign out[2624] = layer_0[11863]; 
    assign out[2625] = ~(layer_0[1480] ^ layer_0[3790]); 
    assign out[2626] = ~layer_0[11368]; 
    assign out[2627] = ~(layer_0[10198] | layer_0[11310]); 
    assign out[2628] = layer_0[7394] & ~layer_0[9947]; 
    assign out[2629] = ~(layer_0[7340] ^ layer_0[10547]); 
    assign out[2630] = ~(layer_0[9564] ^ layer_0[6459]); 
    assign out[2631] = layer_0[2887] ^ layer_0[4864]; 
    assign out[2632] = layer_0[6163] & layer_0[2232]; 
    assign out[2633] = ~(layer_0[6278] ^ layer_0[3702]); 
    assign out[2634] = ~(layer_0[7899] ^ layer_0[11749]); 
    assign out[2635] = layer_0[2673] ^ layer_0[1712]; 
    assign out[2636] = layer_0[1360] ^ layer_0[2659]; 
    assign out[2637] = ~(layer_0[6413] | layer_0[3819]); 
    assign out[2638] = layer_0[3279] ^ layer_0[10687]; 
    assign out[2639] = layer_0[4538] & ~layer_0[29]; 
    assign out[2640] = layer_0[10256]; 
    assign out[2641] = layer_0[7498] & layer_0[2662]; 
    assign out[2642] = ~layer_0[8920] | (layer_0[8920] & layer_0[3626]); 
    assign out[2643] = layer_0[11570]; 
    assign out[2644] = ~(layer_0[11146] ^ layer_0[9585]); 
    assign out[2645] = layer_0[5350] ^ layer_0[502]; 
    assign out[2646] = ~layer_0[6444]; 
    assign out[2647] = ~(layer_0[6294] ^ layer_0[2200]); 
    assign out[2648] = layer_0[4061] ^ layer_0[4186]; 
    assign out[2649] = layer_0[1442] ^ layer_0[10316]; 
    assign out[2650] = layer_0[6814] & layer_0[7136]; 
    assign out[2651] = layer_0[8442] ^ layer_0[11982]; 
    assign out[2652] = layer_0[500] & ~layer_0[3277]; 
    assign out[2653] = layer_0[8742] ^ layer_0[3367]; 
    assign out[2654] = layer_0[11173] & ~layer_0[4745]; 
    assign out[2655] = ~(layer_0[2941] | layer_0[2351]); 
    assign out[2656] = ~layer_0[1395] | (layer_0[2531] & layer_0[1395]); 
    assign out[2657] = layer_0[3450] & ~layer_0[1098]; 
    assign out[2658] = layer_0[2999] ^ layer_0[5581]; 
    assign out[2659] = layer_0[7309] ^ layer_0[10572]; 
    assign out[2660] = layer_0[9313] & ~layer_0[6260]; 
    assign out[2661] = ~(layer_0[11762] ^ layer_0[365]); 
    assign out[2662] = layer_0[104] & ~layer_0[6235]; 
    assign out[2663] = ~layer_0[10095]; 
    assign out[2664] = ~(layer_0[116] ^ layer_0[6406]); 
    assign out[2665] = layer_0[3331] ^ layer_0[3291]; 
    assign out[2666] = layer_0[11995] ^ layer_0[2723]; 
    assign out[2667] = layer_0[3661] & layer_0[10980]; 
    assign out[2668] = layer_0[9144] & ~layer_0[10390]; 
    assign out[2669] = ~(layer_0[9790] ^ layer_0[11149]); 
    assign out[2670] = layer_0[10502] ^ layer_0[1155]; 
    assign out[2671] = layer_0[6120]; 
    assign out[2672] = ~(layer_0[5466] ^ layer_0[3700]); 
    assign out[2673] = ~(layer_0[6363] ^ layer_0[4910]); 
    assign out[2674] = layer_0[11686] ^ layer_0[5411]; 
    assign out[2675] = layer_0[63] ^ layer_0[10247]; 
    assign out[2676] = layer_0[3581] ^ layer_0[6002]; 
    assign out[2677] = ~(layer_0[590] ^ layer_0[2144]); 
    assign out[2678] = ~layer_0[7259]; 
    assign out[2679] = ~layer_0[10704] | (layer_0[10704] & layer_0[4907]); 
    assign out[2680] = layer_0[7597] & layer_0[10250]; 
    assign out[2681] = layer_0[496] & ~layer_0[490]; 
    assign out[2682] = layer_0[10818] & layer_0[7818]; 
    assign out[2683] = ~(layer_0[11152] ^ layer_0[1010]); 
    assign out[2684] = layer_0[6345] ^ layer_0[4152]; 
    assign out[2685] = layer_0[11412] ^ layer_0[5729]; 
    assign out[2686] = layer_0[11799] & ~layer_0[7625]; 
    assign out[2687] = layer_0[1416] ^ layer_0[7784]; 
    assign out[2688] = layer_0[4476] | layer_0[9440]; 
    assign out[2689] = layer_0[6638] ^ layer_0[3048]; 
    assign out[2690] = layer_0[4190]; 
    assign out[2691] = ~(layer_0[151] | layer_0[240]); 
    assign out[2692] = layer_0[3981] ^ layer_0[1589]; 
    assign out[2693] = layer_0[8240] | layer_0[8851]; 
    assign out[2694] = layer_0[9784]; 
    assign out[2695] = layer_0[8208] & layer_0[5001]; 
    assign out[2696] = ~(layer_0[2110] & layer_0[5397]); 
    assign out[2697] = ~(layer_0[10163] & layer_0[11376]); 
    assign out[2698] = layer_0[6072] | layer_0[3547]; 
    assign out[2699] = ~layer_0[1133]; 
    assign out[2700] = ~layer_0[9515] | (layer_0[1827] & layer_0[9515]); 
    assign out[2701] = ~(layer_0[1038] ^ layer_0[1313]); 
    assign out[2702] = ~layer_0[6685] | (layer_0[1742] & layer_0[6685]); 
    assign out[2703] = ~layer_0[3946] | (layer_0[3946] & layer_0[6428]); 
    assign out[2704] = layer_0[9275] ^ layer_0[3252]; 
    assign out[2705] = ~(layer_0[1320] & layer_0[1638]); 
    assign out[2706] = layer_0[2651] & ~layer_0[6670]; 
    assign out[2707] = layer_0[9174] & ~layer_0[3133]; 
    assign out[2708] = ~(layer_0[3470] ^ layer_0[11010]); 
    assign out[2709] = ~(layer_0[9117] ^ layer_0[8258]); 
    assign out[2710] = layer_0[7632] & layer_0[4124]; 
    assign out[2711] = ~(layer_0[5547] ^ layer_0[7056]); 
    assign out[2712] = ~(layer_0[5199] ^ layer_0[8508]); 
    assign out[2713] = layer_0[55] & layer_0[4368]; 
    assign out[2714] = layer_0[6503] & ~layer_0[5415]; 
    assign out[2715] = layer_0[3107] ^ layer_0[9042]; 
    assign out[2716] = layer_0[626] ^ layer_0[6927]; 
    assign out[2717] = ~layer_0[6863]; 
    assign out[2718] = layer_0[5779] & ~layer_0[1292]; 
    assign out[2719] = layer_0[4983] ^ layer_0[9082]; 
    assign out[2720] = layer_0[6262] | layer_0[689]; 
    assign out[2721] = ~(layer_0[3553] ^ layer_0[8688]); 
    assign out[2722] = layer_0[10515] ^ layer_0[6830]; 
    assign out[2723] = ~(layer_0[3436] | layer_0[4645]); 
    assign out[2724] = ~(layer_0[11115] | layer_0[3470]); 
    assign out[2725] = layer_0[149] & ~layer_0[2522]; 
    assign out[2726] = ~(layer_0[6615] ^ layer_0[10887]); 
    assign out[2727] = layer_0[10389]; 
    assign out[2728] = layer_0[5266] & layer_0[10657]; 
    assign out[2729] = ~(layer_0[9980] | layer_0[6431]); 
    assign out[2730] = ~(layer_0[3053] ^ layer_0[1493]); 
    assign out[2731] = ~(layer_0[9540] ^ layer_0[4552]); 
    assign out[2732] = ~layer_0[11891] | (layer_0[11891] & layer_0[5796]); 
    assign out[2733] = ~(layer_0[8106] ^ layer_0[2309]); 
    assign out[2734] = ~layer_0[9115] | (layer_0[7729] & layer_0[9115]); 
    assign out[2735] = layer_0[4070] ^ layer_0[7374]; 
    assign out[2736] = ~layer_0[4536] | (layer_0[3848] & layer_0[4536]); 
    assign out[2737] = layer_0[6725] ^ layer_0[705]; 
    assign out[2738] = layer_0[4481] & ~layer_0[2733]; 
    assign out[2739] = layer_0[2793] & layer_0[8846]; 
    assign out[2740] = ~(layer_0[2682] ^ layer_0[3084]); 
    assign out[2741] = layer_0[7570]; 
    assign out[2742] = layer_0[931] & layer_0[3528]; 
    assign out[2743] = ~(layer_0[9003] | layer_0[7515]); 
    assign out[2744] = layer_0[8150] & layer_0[9535]; 
    assign out[2745] = layer_0[11926] ^ layer_0[315]; 
    assign out[2746] = ~layer_0[1946] | (layer_0[1946] & layer_0[10747]); 
    assign out[2747] = ~layer_0[7707] | (layer_0[10482] & layer_0[7707]); 
    assign out[2748] = ~(layer_0[8299] ^ layer_0[4534]); 
    assign out[2749] = ~layer_0[5448]; 
    assign out[2750] = ~layer_0[9573]; 
    assign out[2751] = layer_0[3597] & ~layer_0[8485]; 
    assign out[2752] = layer_0[4216] ^ layer_0[7291]; 
    assign out[2753] = ~layer_0[11295]; 
    assign out[2754] = layer_0[1182]; 
    assign out[2755] = ~(layer_0[11670] ^ layer_0[4698]); 
    assign out[2756] = layer_0[1751]; 
    assign out[2757] = layer_0[7343] & ~layer_0[8805]; 
    assign out[2758] = ~layer_0[5365]; 
    assign out[2759] = ~(layer_0[2166] ^ layer_0[7069]); 
    assign out[2760] = ~(layer_0[5925] & layer_0[8879]); 
    assign out[2761] = layer_0[5755] ^ layer_0[8946]; 
    assign out[2762] = ~(layer_0[3656] & layer_0[7839]); 
    assign out[2763] = layer_0[566] & ~layer_0[5228]; 
    assign out[2764] = layer_0[3466] ^ layer_0[10942]; 
    assign out[2765] = layer_0[3097] ^ layer_0[312]; 
    assign out[2766] = ~(layer_0[11033] | layer_0[11253]); 
    assign out[2767] = ~layer_0[6477] | (layer_0[6477] & layer_0[7574]); 
    assign out[2768] = layer_0[3933] ^ layer_0[2256]; 
    assign out[2769] = ~layer_0[11345] | (layer_0[11345] & layer_0[10212]); 
    assign out[2770] = layer_0[7580] & ~layer_0[3994]; 
    assign out[2771] = ~layer_0[2685] | (layer_0[4478] & layer_0[2685]); 
    assign out[2772] = layer_0[6739] ^ layer_0[1470]; 
    assign out[2773] = layer_0[576] ^ layer_0[1572]; 
    assign out[2774] = ~(layer_0[5670] ^ layer_0[8032]); 
    assign out[2775] = layer_0[10898] ^ layer_0[4721]; 
    assign out[2776] = layer_0[4500]; 
    assign out[2777] = layer_0[6662] ^ layer_0[7257]; 
    assign out[2778] = layer_0[7589] ^ layer_0[7120]; 
    assign out[2779] = layer_0[554] & layer_0[6448]; 
    assign out[2780] = layer_0[10488] ^ layer_0[7876]; 
    assign out[2781] = ~(layer_0[4928] ^ layer_0[10746]); 
    assign out[2782] = ~layer_0[6703]; 
    assign out[2783] = layer_0[8126]; 
    assign out[2784] = layer_0[667] ^ layer_0[6455]; 
    assign out[2785] = layer_0[7241] ^ layer_0[2849]; 
    assign out[2786] = layer_0[11198] & ~layer_0[8720]; 
    assign out[2787] = layer_0[8026] & ~layer_0[8674]; 
    assign out[2788] = layer_0[8511] ^ layer_0[2833]; 
    assign out[2789] = ~(layer_0[8122] ^ layer_0[2758]); 
    assign out[2790] = ~layer_0[9379] | (layer_0[9379] & layer_0[6347]); 
    assign out[2791] = ~layer_0[5549] | (layer_0[5549] & layer_0[10274]); 
    assign out[2792] = layer_0[1635] | layer_0[4050]; 
    assign out[2793] = ~(layer_0[3134] ^ layer_0[9314]); 
    assign out[2794] = ~(layer_0[2549] ^ layer_0[9146]); 
    assign out[2795] = ~(layer_0[1548] ^ layer_0[10111]); 
    assign out[2796] = ~layer_0[11661] | (layer_0[4572] & layer_0[11661]); 
    assign out[2797] = layer_0[2628] ^ layer_0[11949]; 
    assign out[2798] = layer_0[9814] ^ layer_0[2179]; 
    assign out[2799] = ~(layer_0[3825] ^ layer_0[3906]); 
    assign out[2800] = layer_0[8967] ^ layer_0[7313]; 
    assign out[2801] = ~(layer_0[8691] ^ layer_0[328]); 
    assign out[2802] = layer_0[8900]; 
    assign out[2803] = layer_0[9371] ^ layer_0[4185]; 
    assign out[2804] = ~(layer_0[8326] ^ layer_0[7539]); 
    assign out[2805] = ~(layer_0[11754] & layer_0[2581]); 
    assign out[2806] = layer_0[9859] ^ layer_0[11468]; 
    assign out[2807] = layer_0[9583] | layer_0[1864]; 
    assign out[2808] = layer_0[3781] ^ layer_0[11569]; 
    assign out[2809] = ~(layer_0[494] ^ layer_0[9027]); 
    assign out[2810] = layer_0[349]; 
    assign out[2811] = layer_0[9139] & ~layer_0[228]; 
    assign out[2812] = ~(layer_0[8305] ^ layer_0[9472]); 
    assign out[2813] = ~(layer_0[9107] ^ layer_0[11045]); 
    assign out[2814] = ~(layer_0[651] | layer_0[3296]); 
    assign out[2815] = layer_0[8780] ^ layer_0[7582]; 
    assign out[2816] = ~(layer_0[5947] ^ layer_0[7892]); 
    assign out[2817] = layer_0[7577] & layer_0[7789]; 
    assign out[2818] = ~(layer_0[5019] ^ layer_0[5981]); 
    assign out[2819] = ~layer_0[5409] | (layer_0[9884] & layer_0[5409]); 
    assign out[2820] = ~layer_0[4566]; 
    assign out[2821] = ~layer_0[10127] | (layer_0[10653] & layer_0[10127]); 
    assign out[2822] = ~(layer_0[1078] ^ layer_0[9419]); 
    assign out[2823] = layer_0[8196] | layer_0[4554]; 
    assign out[2824] = ~(layer_0[2726] | layer_0[6708]); 
    assign out[2825] = layer_0[6562] ^ layer_0[8539]; 
    assign out[2826] = ~(layer_0[5015] ^ layer_0[2345]); 
    assign out[2827] = ~layer_0[3087]; 
    assign out[2828] = layer_0[2360] & layer_0[2201]; 
    assign out[2829] = ~(layer_0[4711] ^ layer_0[4939]); 
    assign out[2830] = layer_0[565] ^ layer_0[8687]; 
    assign out[2831] = ~(layer_0[9433] ^ layer_0[9349]); 
    assign out[2832] = ~layer_0[1344]; 
    assign out[2833] = layer_0[9344]; 
    assign out[2834] = ~(layer_0[4116] ^ layer_0[4240]); 
    assign out[2835] = ~(layer_0[6083] ^ layer_0[10099]); 
    assign out[2836] = ~(layer_0[48] ^ layer_0[8544]); 
    assign out[2837] = ~(layer_0[5014] ^ layer_0[4431]); 
    assign out[2838] = layer_0[11714] ^ layer_0[5209]; 
    assign out[2839] = ~(layer_0[5356] & layer_0[1998]); 
    assign out[2840] = layer_0[5479]; 
    assign out[2841] = ~(layer_0[5907] ^ layer_0[9572]); 
    assign out[2842] = layer_0[2542] ^ layer_0[8860]; 
    assign out[2843] = layer_0[7946] ^ layer_0[5846]; 
    assign out[2844] = ~layer_0[4775]; 
    assign out[2845] = ~layer_0[7546] | (layer_0[7546] & layer_0[5568]); 
    assign out[2846] = layer_0[8704]; 
    assign out[2847] = ~layer_0[1025]; 
    assign out[2848] = layer_0[7428] ^ layer_0[10392]; 
    assign out[2849] = ~layer_0[8012] | (layer_0[8012] & layer_0[5414]); 
    assign out[2850] = layer_0[11943] & layer_0[9010]; 
    assign out[2851] = ~(layer_0[2395] ^ layer_0[2569]); 
    assign out[2852] = ~layer_0[2738] | (layer_0[2738] & layer_0[7779]); 
    assign out[2853] = ~(layer_0[5999] ^ layer_0[374]); 
    assign out[2854] = layer_0[572] | layer_0[646]; 
    assign out[2855] = ~layer_0[10026]; 
    assign out[2856] = ~layer_0[11817] | (layer_0[133] & layer_0[11817]); 
    assign out[2857] = ~(layer_0[11636] ^ layer_0[8365]); 
    assign out[2858] = ~(layer_0[980] ^ layer_0[8605]); 
    assign out[2859] = layer_0[1765] & ~layer_0[2171]; 
    assign out[2860] = ~(layer_0[9460] ^ layer_0[6241]); 
    assign out[2861] = layer_0[646] ^ layer_0[2886]; 
    assign out[2862] = ~layer_0[3777]; 
    assign out[2863] = layer_0[8735]; 
    assign out[2864] = layer_0[1233] ^ layer_0[10547]; 
    assign out[2865] = ~(layer_0[7967] ^ layer_0[7081]); 
    assign out[2866] = ~(layer_0[6520] ^ layer_0[10440]); 
    assign out[2867] = layer_0[5044] ^ layer_0[4208]; 
    assign out[2868] = ~layer_0[13]; 
    assign out[2869] = layer_0[11401] & ~layer_0[7476]; 
    assign out[2870] = ~(layer_0[7481] ^ layer_0[10709]); 
    assign out[2871] = layer_0[11426] ^ layer_0[5255]; 
    assign out[2872] = ~(layer_0[3018] ^ layer_0[7210]); 
    assign out[2873] = layer_0[8634] ^ layer_0[336]; 
    assign out[2874] = ~(layer_0[9800] ^ layer_0[2623]); 
    assign out[2875] = ~layer_0[8063] | (layer_0[8063] & layer_0[6911]); 
    assign out[2876] = ~(layer_0[7373] ^ layer_0[414]); 
    assign out[2877] = ~layer_0[3444]; 
    assign out[2878] = ~(layer_0[4181] ^ layer_0[4881]); 
    assign out[2879] = ~layer_0[1760] | (layer_0[10126] & layer_0[1760]); 
    assign out[2880] = ~(layer_0[7617] ^ layer_0[6960]); 
    assign out[2881] = ~layer_0[3087] | (layer_0[3087] & layer_0[734]); 
    assign out[2882] = layer_0[11441] & ~layer_0[3731]; 
    assign out[2883] = ~(layer_0[10494] ^ layer_0[10439]); 
    assign out[2884] = layer_0[6313] ^ layer_0[11809]; 
    assign out[2885] = ~(layer_0[9238] ^ layer_0[6211]); 
    assign out[2886] = layer_0[8973] & ~layer_0[5795]; 
    assign out[2887] = layer_0[2462] ^ layer_0[2061]; 
    assign out[2888] = ~layer_0[3982]; 
    assign out[2889] = layer_0[6282] ^ layer_0[10257]; 
    assign out[2890] = layer_0[7752] ^ layer_0[9271]; 
    assign out[2891] = ~(layer_0[624] ^ layer_0[9366]); 
    assign out[2892] = ~(layer_0[2711] ^ layer_0[5804]); 
    assign out[2893] = ~(layer_0[4792] ^ layer_0[9594]); 
    assign out[2894] = layer_0[4450]; 
    assign out[2895] = layer_0[11150]; 
    assign out[2896] = layer_0[6193] ^ layer_0[2712]; 
    assign out[2897] = layer_0[6305]; 
    assign out[2898] = layer_0[8233] ^ layer_0[1466]; 
    assign out[2899] = ~(layer_0[11299] ^ layer_0[6582]); 
    assign out[2900] = ~layer_0[8024] | (layer_0[8024] & layer_0[11900]); 
    assign out[2901] = ~layer_0[7014]; 
    assign out[2902] = ~(layer_0[9545] | layer_0[8719]); 
    assign out[2903] = layer_0[10316] ^ layer_0[11639]; 
    assign out[2904] = ~layer_0[9617]; 
    assign out[2905] = layer_0[10380] ^ layer_0[8773]; 
    assign out[2906] = layer_0[4809]; 
    assign out[2907] = layer_0[4719] & ~layer_0[3829]; 
    assign out[2908] = layer_0[6825] | layer_0[11548]; 
    assign out[2909] = ~(layer_0[6421] ^ layer_0[4844]); 
    assign out[2910] = ~(layer_0[4253] ^ layer_0[9358]); 
    assign out[2911] = ~(layer_0[2006] ^ layer_0[10268]); 
    assign out[2912] = ~(layer_0[8167] ^ layer_0[8686]); 
    assign out[2913] = ~(layer_0[5212] ^ layer_0[4146]); 
    assign out[2914] = layer_0[9322]; 
    assign out[2915] = layer_0[6567] ^ layer_0[11649]; 
    assign out[2916] = ~(layer_0[10056] ^ layer_0[9867]); 
    assign out[2917] = layer_0[10699] & ~layer_0[769]; 
    assign out[2918] = layer_0[165] & layer_0[10602]; 
    assign out[2919] = ~layer_0[6762]; 
    assign out[2920] = ~(layer_0[10640] | layer_0[2593]); 
    assign out[2921] = layer_0[418] & ~layer_0[9526]; 
    assign out[2922] = layer_0[4339] ^ layer_0[6515]; 
    assign out[2923] = layer_0[9201] ^ layer_0[3373]; 
    assign out[2924] = layer_0[11104] ^ layer_0[4307]; 
    assign out[2925] = ~(layer_0[4199] ^ layer_0[5284]); 
    assign out[2926] = layer_0[9402] & ~layer_0[997]; 
    assign out[2927] = layer_0[7296] | layer_0[229]; 
    assign out[2928] = layer_0[8204] & ~layer_0[6573]; 
    assign out[2929] = layer_0[5843] ^ layer_0[3802]; 
    assign out[2930] = layer_0[11928] ^ layer_0[367]; 
    assign out[2931] = layer_0[2360] ^ layer_0[10782]; 
    assign out[2932] = layer_0[7593] & ~layer_0[4389]; 
    assign out[2933] = ~(layer_0[2629] ^ layer_0[1185]); 
    assign out[2934] = ~(layer_0[9410] & layer_0[11907]); 
    assign out[2935] = ~layer_0[10687] | (layer_0[11294] & layer_0[10687]); 
    assign out[2936] = ~layer_0[3334]; 
    assign out[2937] = ~layer_0[7694]; 
    assign out[2938] = ~(layer_0[6917] ^ layer_0[9740]); 
    assign out[2939] = layer_0[4180] ^ layer_0[8554]; 
    assign out[2940] = layer_0[6105] & ~layer_0[345]; 
    assign out[2941] = layer_0[5470] ^ layer_0[6900]; 
    assign out[2942] = layer_0[10145] & layer_0[5718]; 
    assign out[2943] = ~(layer_0[10334] ^ layer_0[5003]); 
    assign out[2944] = layer_0[11767] ^ layer_0[4659]; 
    assign out[2945] = ~layer_0[7128] | (layer_0[7128] & layer_0[4258]); 
    assign out[2946] = ~(layer_0[6121] & layer_0[8393]); 
    assign out[2947] = ~(layer_0[2193] ^ layer_0[6783]); 
    assign out[2948] = layer_0[2481] & ~layer_0[6946]; 
    assign out[2949] = layer_0[5224] ^ layer_0[3032]; 
    assign out[2950] = layer_0[6202] & layer_0[11666]; 
    assign out[2951] = layer_0[4063] | layer_0[5860]; 
    assign out[2952] = layer_0[1573] ^ layer_0[2586]; 
    assign out[2953] = layer_0[1356]; 
    assign out[2954] = layer_0[640] ^ layer_0[10957]; 
    assign out[2955] = layer_0[7673] & layer_0[11628]; 
    assign out[2956] = ~(layer_0[551] ^ layer_0[7017]); 
    assign out[2957] = ~(layer_0[9380] ^ layer_0[10683]); 
    assign out[2958] = layer_0[5635] ^ layer_0[6380]; 
    assign out[2959] = layer_0[9509] ^ layer_0[9290]; 
    assign out[2960] = ~(layer_0[7112] ^ layer_0[3293]); 
    assign out[2961] = ~layer_0[7375]; 
    assign out[2962] = layer_0[8082] ^ layer_0[5677]; 
    assign out[2963] = layer_0[739]; 
    assign out[2964] = layer_0[9315] ^ layer_0[5753]; 
    assign out[2965] = ~(layer_0[4217] & layer_0[2638]); 
    assign out[2966] = layer_0[6647] ^ layer_0[2716]; 
    assign out[2967] = ~layer_0[7443] | (layer_0[4667] & layer_0[7443]); 
    assign out[2968] = ~(layer_0[2591] ^ layer_0[2303]); 
    assign out[2969] = ~(layer_0[1346] ^ layer_0[11492]); 
    assign out[2970] = ~layer_0[5936]; 
    assign out[2971] = ~(layer_0[8523] ^ layer_0[10714]); 
    assign out[2972] = ~layer_0[4602]; 
    assign out[2973] = ~layer_0[10560]; 
    assign out[2974] = layer_0[3858] & layer_0[5910]; 
    assign out[2975] = layer_0[5026] ^ layer_0[11956]; 
    assign out[2976] = ~(layer_0[9053] | layer_0[8125]); 
    assign out[2977] = ~(layer_0[11402] ^ layer_0[6999]); 
    assign out[2978] = layer_0[8832]; 
    assign out[2979] = layer_0[7073] ^ layer_0[3704]; 
    assign out[2980] = ~(layer_0[241] ^ layer_0[6189]); 
    assign out[2981] = layer_0[7337] & layer_0[4796]; 
    assign out[2982] = ~layer_0[11181] | (layer_0[4816] & layer_0[11181]); 
    assign out[2983] = ~(layer_0[9365] | layer_0[10369]); 
    assign out[2984] = ~layer_0[8890]; 
    assign out[2985] = layer_0[8929] ^ layer_0[3583]; 
    assign out[2986] = ~(layer_0[3720] & layer_0[6485]); 
    assign out[2987] = layer_0[6124] ^ layer_0[6152]; 
    assign out[2988] = ~(layer_0[11864] | layer_0[6144]); 
    assign out[2989] = layer_0[1256] ^ layer_0[11502]; 
    assign out[2990] = layer_0[309] | layer_0[4673]; 
    assign out[2991] = layer_0[4898] ^ layer_0[973]; 
    assign out[2992] = layer_0[2100]; 
    assign out[2993] = ~layer_0[5959]; 
    assign out[2994] = layer_0[3958] ^ layer_0[10116]; 
    assign out[2995] = ~(layer_0[5765] ^ layer_0[6744]); 
    assign out[2996] = ~layer_0[239] | (layer_0[239] & layer_0[5297]); 
    assign out[2997] = layer_0[7871]; 
    assign out[2998] = layer_0[1722] ^ layer_0[8029]; 
    assign out[2999] = layer_0[5731] ^ layer_0[4741]; 
    assign out[3000] = ~(layer_0[6565] ^ layer_0[6611]); 
    assign out[3001] = layer_0[10181]; 
    assign out[3002] = layer_0[8311] ^ layer_0[3283]; 
    assign out[3003] = layer_0[96] ^ layer_0[7691]; 
    assign out[3004] = layer_0[87] ^ layer_0[9828]; 
    assign out[3005] = layer_0[50] ^ layer_0[4223]; 
    assign out[3006] = ~layer_0[11055] | (layer_0[9930] & layer_0[11055]); 
    assign out[3007] = ~(layer_0[5840] ^ layer_0[4540]); 
    assign out[3008] = ~(layer_0[11372] ^ layer_0[5698]); 
    assign out[3009] = layer_0[1944] & ~layer_0[9719]; 
    assign out[3010] = ~layer_0[9380] | (layer_0[9380] & layer_0[4575]); 
    assign out[3011] = ~layer_0[2701]; 
    assign out[3012] = ~(layer_0[9320] ^ layer_0[534]); 
    assign out[3013] = layer_0[7920]; 
    assign out[3014] = layer_0[7417] & ~layer_0[8703]; 
    assign out[3015] = layer_0[11499]; 
    assign out[3016] = ~layer_0[11308] | (layer_0[11308] & layer_0[9105]); 
    assign out[3017] = ~(layer_0[3689] ^ layer_0[11572]); 
    assign out[3018] = layer_0[3784] & ~layer_0[5577]; 
    assign out[3019] = layer_0[7552] | layer_0[3401]; 
    assign out[3020] = ~(layer_0[6228] | layer_0[3554]); 
    assign out[3021] = ~layer_0[5488] | (layer_0[5488] & layer_0[5625]); 
    assign out[3022] = ~layer_0[2615] | (layer_0[2059] & layer_0[2615]); 
    assign out[3023] = layer_0[1117] ^ layer_0[511]; 
    assign out[3024] = ~(layer_0[11871] ^ layer_0[5725]); 
    assign out[3025] = ~(layer_0[4559] ^ layer_0[7012]); 
    assign out[3026] = layer_0[11524] & ~layer_0[7348]; 
    assign out[3027] = ~(layer_0[4922] & layer_0[2782]); 
    assign out[3028] = ~(layer_0[1532] | layer_0[6079]); 
    assign out[3029] = layer_0[4523] & ~layer_0[4596]; 
    assign out[3030] = layer_0[1894]; 
    assign out[3031] = ~(layer_0[8021] & layer_0[5803]); 
    assign out[3032] = layer_0[5169]; 
    assign out[3033] = layer_0[4077] & layer_0[10715]; 
    assign out[3034] = layer_0[7127] ^ layer_0[11217]; 
    assign out[3035] = ~layer_0[6568]; 
    assign out[3036] = layer_0[3892]; 
    assign out[3037] = layer_0[7359] ^ layer_0[11165]; 
    assign out[3038] = ~(layer_0[5204] ^ layer_0[9325]); 
    assign out[3039] = ~(layer_0[1748] ^ layer_0[2565]); 
    assign out[3040] = layer_0[8168] & ~layer_0[7387]; 
    assign out[3041] = ~layer_0[8608]; 
    assign out[3042] = layer_0[3785] & layer_0[6883]; 
    assign out[3043] = layer_0[11778] & ~layer_0[2227]; 
    assign out[3044] = layer_0[10624] ^ layer_0[6123]; 
    assign out[3045] = ~(layer_0[9742] | layer_0[933]); 
    assign out[3046] = ~layer_0[4072]; 
    assign out[3047] = layer_0[2827] & ~layer_0[421]; 
    assign out[3048] = layer_0[2062] ^ layer_0[8514]; 
    assign out[3049] = layer_0[373] ^ layer_0[10712]; 
    assign out[3050] = layer_0[860] & ~layer_0[1749]; 
    assign out[3051] = layer_0[2656] & ~layer_0[7832]; 
    assign out[3052] = layer_0[7663] & ~layer_0[3877]; 
    assign out[3053] = ~layer_0[4977] | (layer_0[4977] & layer_0[2894]); 
    assign out[3054] = layer_0[7985] ^ layer_0[2567]; 
    assign out[3055] = layer_0[9166] ^ layer_0[8371]; 
    assign out[3056] = layer_0[5160]; 
    assign out[3057] = ~layer_0[225]; 
    assign out[3058] = ~(layer_0[7322] ^ layer_0[9847]); 
    assign out[3059] = ~(layer_0[1200] ^ layer_0[6068]); 
    assign out[3060] = layer_0[2902] | layer_0[10503]; 
    assign out[3061] = layer_0[9925] ^ layer_0[6418]; 
    assign out[3062] = layer_0[5418] & ~layer_0[6025]; 
    assign out[3063] = ~(layer_0[4447] ^ layer_0[11163]); 
    assign out[3064] = layer_0[727] & ~layer_0[8820]; 
    assign out[3065] = ~(layer_0[9310] ^ layer_0[4578]); 
    assign out[3066] = layer_0[8646] & ~layer_0[10701]; 
    assign out[3067] = layer_0[9835] & ~layer_0[2695]; 
    assign out[3068] = ~(layer_0[11071] ^ layer_0[7388]); 
    assign out[3069] = ~(layer_0[10550] ^ layer_0[3990]); 
    assign out[3070] = ~(layer_0[5364] ^ layer_0[11285]); 
    assign out[3071] = ~(layer_0[5403] ^ layer_0[9345]); 
    assign out[3072] = ~(layer_0[5456] | layer_0[6835]); 
    assign out[3073] = layer_0[1049] & ~layer_0[2425]; 
    assign out[3074] = ~(layer_0[7485] ^ layer_0[2591]); 
    assign out[3075] = ~(layer_0[11383] ^ layer_0[7545]); 
    assign out[3076] = layer_0[10335] & ~layer_0[6558]; 
    assign out[3077] = ~(layer_0[1939] | layer_0[7003]); 
    assign out[3078] = layer_0[1421] & ~layer_0[7129]; 
    assign out[3079] = layer_0[11852] ^ layer_0[11185]; 
    assign out[3080] = ~(layer_0[1216] ^ layer_0[1481]); 
    assign out[3081] = ~(layer_0[5136] ^ layer_0[423]); 
    assign out[3082] = layer_0[7175] ^ layer_0[100]; 
    assign out[3083] = layer_0[426] & layer_0[11112]; 
    assign out[3084] = ~(layer_0[2730] ^ layer_0[3272]); 
    assign out[3085] = ~(layer_0[8259] ^ layer_0[1163]); 
    assign out[3086] = layer_0[2749] & ~layer_0[6527]; 
    assign out[3087] = ~layer_0[3932] | (layer_0[7761] & layer_0[3932]); 
    assign out[3088] = layer_0[5509] ^ layer_0[4931]; 
    assign out[3089] = ~layer_0[9688]; 
    assign out[3090] = ~(layer_0[552] ^ layer_0[6252]); 
    assign out[3091] = ~(layer_0[7918] | layer_0[6898]); 
    assign out[3092] = layer_0[552] ^ layer_0[6712]; 
    assign out[3093] = layer_0[10050] ^ layer_0[1581]; 
    assign out[3094] = ~layer_0[4035]; 
    assign out[3095] = ~(layer_0[863] ^ layer_0[10129]); 
    assign out[3096] = layer_0[11608] ^ layer_0[2041]; 
    assign out[3097] = ~(layer_0[8121] | layer_0[7200]); 
    assign out[3098] = layer_0[7115] & layer_0[11531]; 
    assign out[3099] = ~(layer_0[535] ^ layer_0[1465]); 
    assign out[3100] = ~(layer_0[3840] ^ layer_0[1102]); 
    assign out[3101] = ~layer_0[5406]; 
    assign out[3102] = layer_0[2176]; 
    assign out[3103] = ~(layer_0[2992] ^ layer_0[4996]); 
    assign out[3104] = ~(layer_0[1453] ^ layer_0[8306]); 
    assign out[3105] = ~(layer_0[8397] ^ layer_0[11623]); 
    assign out[3106] = layer_0[7563]; 
    assign out[3107] = layer_0[1419] & ~layer_0[6115]; 
    assign out[3108] = layer_0[4505] ^ layer_0[3608]; 
    assign out[3109] = layer_0[9494] & layer_0[10608]; 
    assign out[3110] = layer_0[6424] ^ layer_0[4096]; 
    assign out[3111] = ~(layer_0[10492] ^ layer_0[6704]); 
    assign out[3112] = layer_0[9751] & layer_0[9754]; 
    assign out[3113] = layer_0[2291] ^ layer_0[6251]; 
    assign out[3114] = layer_0[7403] ^ layer_0[8383]; 
    assign out[3115] = layer_0[2225] ^ layer_0[1110]; 
    assign out[3116] = layer_0[7578] ^ layer_0[10352]; 
    assign out[3117] = layer_0[3162] ^ layer_0[8134]; 
    assign out[3118] = layer_0[2347] & layer_0[5412]; 
    assign out[3119] = ~(layer_0[3766] ^ layer_0[5676]); 
    assign out[3120] = layer_0[627] ^ layer_0[574]; 
    assign out[3121] = ~(layer_0[3244] ^ layer_0[10014]); 
    assign out[3122] = ~layer_0[1966] | (layer_0[528] & layer_0[1966]); 
    assign out[3123] = layer_0[10581] ^ layer_0[11291]; 
    assign out[3124] = layer_0[10419]; 
    assign out[3125] = ~layer_0[4678]; 
    assign out[3126] = layer_0[9075]; 
    assign out[3127] = layer_0[4040] ^ layer_0[9220]; 
    assign out[3128] = layer_0[4963] & ~layer_0[11615]; 
    assign out[3129] = ~(layer_0[5374] ^ layer_0[11438]); 
    assign out[3130] = ~layer_0[2854] | (layer_0[2854] & layer_0[11620]); 
    assign out[3131] = layer_0[638] | layer_0[6607]; 
    assign out[3132] = ~(layer_0[7385] ^ layer_0[11770]); 
    assign out[3133] = ~(layer_0[4022] ^ layer_0[1755]); 
    assign out[3134] = layer_0[7323] & layer_0[9992]; 
    assign out[3135] = ~(layer_0[5941] ^ layer_0[11030]); 
    assign out[3136] = layer_0[9394] ^ layer_0[4343]; 
    assign out[3137] = ~(layer_0[6188] ^ layer_0[3975]); 
    assign out[3138] = ~layer_0[11948]; 
    assign out[3139] = ~layer_0[1879]; 
    assign out[3140] = layer_0[8859]; 
    assign out[3141] = ~layer_0[1611]; 
    assign out[3142] = ~(layer_0[4413] | layer_0[10384]); 
    assign out[3143] = layer_0[5582] ^ layer_0[716]; 
    assign out[3144] = ~layer_0[7289] | (layer_0[7289] & layer_0[6598]); 
    assign out[3145] = ~(layer_0[6919] & layer_0[2659]); 
    assign out[3146] = layer_0[966]; 
    assign out[3147] = layer_0[725] & layer_0[1660]; 
    assign out[3148] = layer_0[5863] | layer_0[7310]; 
    assign out[3149] = ~layer_0[3185]; 
    assign out[3150] = ~layer_0[8350]; 
    assign out[3151] = layer_0[1592] ^ layer_0[2558]; 
    assign out[3152] = layer_0[7305] ^ layer_0[2479]; 
    assign out[3153] = layer_0[7713]; 
    assign out[3154] = ~layer_0[11503]; 
    assign out[3155] = ~layer_0[5424] | (layer_0[1677] & layer_0[5424]); 
    assign out[3156] = layer_0[5988] ^ layer_0[7680]; 
    assign out[3157] = layer_0[8512] & layer_0[8971]; 
    assign out[3158] = layer_0[8262] ^ layer_0[11414]; 
    assign out[3159] = ~layer_0[4851]; 
    assign out[3160] = ~(layer_0[3778] ^ layer_0[3177]); 
    assign out[3161] = layer_0[1778]; 
    assign out[3162] = ~(layer_0[11937] ^ layer_0[5982]); 
    assign out[3163] = ~(layer_0[5462] ^ layer_0[4987]); 
    assign out[3164] = ~layer_0[10338]; 
    assign out[3165] = layer_0[8233] ^ layer_0[1027]; 
    assign out[3166] = layer_0[2111] ^ layer_0[404]; 
    assign out[3167] = layer_0[662]; 
    assign out[3168] = layer_0[3396] ^ layer_0[10088]; 
    assign out[3169] = ~(layer_0[10428] ^ layer_0[3438]); 
    assign out[3170] = layer_0[884]; 
    assign out[3171] = ~layer_0[8076]; 
    assign out[3172] = ~(layer_0[9265] & layer_0[2678]); 
    assign out[3173] = layer_0[870] ^ layer_0[1542]; 
    assign out[3174] = ~layer_0[675]; 
    assign out[3175] = layer_0[9722] ^ layer_0[8981]; 
    assign out[3176] = ~layer_0[364] | (layer_0[2881] & layer_0[364]); 
    assign out[3177] = layer_0[6713] ^ layer_0[7469]; 
    assign out[3178] = layer_0[2412]; 
    assign out[3179] = layer_0[9184] ^ layer_0[9751]; 
    assign out[3180] = ~(layer_0[6578] ^ layer_0[6240]); 
    assign out[3181] = ~(layer_0[6470] ^ layer_0[3148]); 
    assign out[3182] = layer_0[8882] & ~layer_0[10219]; 
    assign out[3183] = layer_0[5504]; 
    assign out[3184] = ~(layer_0[5908] ^ layer_0[924]); 
    assign out[3185] = layer_0[9619] ^ layer_0[4759]; 
    assign out[3186] = ~layer_0[9286]; 
    assign out[3187] = ~layer_0[6956] | (layer_0[6956] & layer_0[8426]); 
    assign out[3188] = ~layer_0[8266] | (layer_0[8266] & layer_0[2213]); 
    assign out[3189] = ~(layer_0[8966] ^ layer_0[11561]); 
    assign out[3190] = ~(layer_0[4664] ^ layer_0[3937]); 
    assign out[3191] = ~(layer_0[6589] ^ layer_0[1552]); 
    assign out[3192] = ~(layer_0[2038] ^ layer_0[7149]); 
    assign out[3193] = ~(layer_0[11141] ^ layer_0[10442]); 
    assign out[3194] = layer_0[11819] ^ layer_0[734]; 
    assign out[3195] = ~(layer_0[8728] ^ layer_0[10991]); 
    assign out[3196] = ~(layer_0[9197] ^ layer_0[10779]); 
    assign out[3197] = layer_0[329] ^ layer_0[3140]; 
    assign out[3198] = ~(layer_0[11279] ^ layer_0[4654]); 
    assign out[3199] = layer_0[10147] ^ layer_0[3833]; 
    assign out[3200] = layer_0[8104] ^ layer_0[11508]; 
    assign out[3201] = layer_0[2279] & layer_0[6036]; 
    assign out[3202] = ~(layer_0[6283] ^ layer_0[2487]); 
    assign out[3203] = layer_0[4641] ^ layer_0[10502]; 
    assign out[3204] = layer_0[751] & ~layer_0[8816]; 
    assign out[3205] = ~(layer_0[6677] ^ layer_0[3128]); 
    assign out[3206] = layer_0[9482] & ~layer_0[2088]; 
    assign out[3207] = layer_0[8855] & ~layer_0[5318]; 
    assign out[3208] = ~layer_0[5822]; 
    assign out[3209] = ~(layer_0[1725] ^ layer_0[9442]); 
    assign out[3210] = layer_0[9288] | layer_0[7517]; 
    assign out[3211] = ~(layer_0[3431] ^ layer_0[515]); 
    assign out[3212] = ~layer_0[3480] | (layer_0[4556] & layer_0[3480]); 
    assign out[3213] = ~layer_0[570]; 
    assign out[3214] = ~(layer_0[10663] ^ layer_0[699]); 
    assign out[3215] = layer_0[8532]; 
    assign out[3216] = ~(layer_0[2924] ^ layer_0[3568]); 
    assign out[3217] = ~(layer_0[11676] ^ layer_0[5758]); 
    assign out[3218] = ~(layer_0[2298] | layer_0[1149]); 
    assign out[3219] = layer_0[7584] & layer_0[10812]; 
    assign out[3220] = layer_0[7380] ^ layer_0[1563]; 
    assign out[3221] = layer_0[2819] ^ layer_0[1764]; 
    assign out[3222] = layer_0[2663] ^ layer_0[529]; 
    assign out[3223] = layer_0[4707] & layer_0[9839]; 
    assign out[3224] = layer_0[8489] & ~layer_0[68]; 
    assign out[3225] = layer_0[5523] & ~layer_0[806]; 
    assign out[3226] = layer_0[4688] ^ layer_0[6683]; 
    assign out[3227] = layer_0[7140] ^ layer_0[8308]; 
    assign out[3228] = layer_0[1633] & layer_0[79]; 
    assign out[3229] = layer_0[3878]; 
    assign out[3230] = ~(layer_0[5062] | layer_0[4400]); 
    assign out[3231] = layer_0[1477] ^ layer_0[1862]; 
    assign out[3232] = ~layer_0[10007] | (layer_0[10007] & layer_0[10724]); 
    assign out[3233] = layer_0[10652] ^ layer_0[7312]; 
    assign out[3234] = layer_0[11826]; 
    assign out[3235] = ~(layer_0[2320] ^ layer_0[7127]); 
    assign out[3236] = layer_0[2952] ^ layer_0[858]; 
    assign out[3237] = layer_0[4674] ^ layer_0[6969]; 
    assign out[3238] = layer_0[7638] ^ layer_0[253]; 
    assign out[3239] = layer_0[8466] & layer_0[3482]; 
    assign out[3240] = ~(layer_0[6895] ^ layer_0[3064]); 
    assign out[3241] = layer_0[10841] & layer_0[6984]; 
    assign out[3242] = ~(layer_0[10232] ^ layer_0[4419]); 
    assign out[3243] = ~layer_0[4633] | (layer_0[4633] & layer_0[9864]); 
    assign out[3244] = ~(layer_0[5865] | layer_0[1964]); 
    assign out[3245] = layer_0[10431] & ~layer_0[1053]; 
    assign out[3246] = layer_0[3818]; 
    assign out[3247] = layer_0[3108] ^ layer_0[8377]; 
    assign out[3248] = layer_0[8002] ^ layer_0[1042]; 
    assign out[3249] = ~(layer_0[1358] | layer_0[3]); 
    assign out[3250] = layer_0[4599]; 
    assign out[3251] = ~(layer_0[300] ^ layer_0[9373]); 
    assign out[3252] = ~(layer_0[5072] | layer_0[11750]); 
    assign out[3253] = layer_0[7497] ^ layer_0[563]; 
    assign out[3254] = ~(layer_0[3529] ^ layer_0[10998]); 
    assign out[3255] = layer_0[5227] ^ layer_0[3604]; 
    assign out[3256] = layer_0[729] ^ layer_0[183]; 
    assign out[3257] = layer_0[7678]; 
    assign out[3258] = layer_0[3820] & layer_0[9499]; 
    assign out[3259] = layer_0[706] & ~layer_0[8974]; 
    assign out[3260] = layer_0[10585] ^ layer_0[5569]; 
    assign out[3261] = layer_0[452] & ~layer_0[5068]; 
    assign out[3262] = layer_0[8294]; 
    assign out[3263] = ~layer_0[7702] | (layer_0[7702] & layer_0[9273]); 
    assign out[3264] = ~(layer_0[994] ^ layer_0[8887]); 
    assign out[3265] = layer_0[1145] & ~layer_0[1640]; 
    assign out[3266] = layer_0[736] ^ layer_0[5314]; 
    assign out[3267] = ~(layer_0[7261] | layer_0[996]); 
    assign out[3268] = layer_0[11104] & ~layer_0[11351]; 
    assign out[3269] = layer_0[6433] ^ layer_0[6695]; 
    assign out[3270] = layer_0[8586] ^ layer_0[11489]; 
    assign out[3271] = ~layer_0[1678]; 
    assign out[3272] = layer_0[3416] & layer_0[8172]; 
    assign out[3273] = layer_0[7666] & ~layer_0[2879]; 
    assign out[3274] = layer_0[5629] ^ layer_0[8455]; 
    assign out[3275] = ~(layer_0[9283] | layer_0[3750]); 
    assign out[3276] = ~(layer_0[1043] ^ layer_0[7092]); 
    assign out[3277] = ~(layer_0[3007] ^ layer_0[4565]); 
    assign out[3278] = layer_0[7311] ^ layer_0[10089]; 
    assign out[3279] = layer_0[10592] & ~layer_0[49]; 
    assign out[3280] = ~(layer_0[9087] ^ layer_0[10812]); 
    assign out[3281] = ~layer_0[9707] | (layer_0[9707] & layer_0[3538]); 
    assign out[3282] = layer_0[1021]; 
    assign out[3283] = layer_0[9114] & layer_0[5264]; 
    assign out[3284] = ~layer_0[2282]; 
    assign out[3285] = layer_0[5532] ^ layer_0[902]; 
    assign out[3286] = layer_0[8456] & ~layer_0[4824]; 
    assign out[3287] = ~(layer_0[2106] ^ layer_0[2275]); 
    assign out[3288] = layer_0[5334] & ~layer_0[10185]; 
    assign out[3289] = layer_0[1] ^ layer_0[9022]; 
    assign out[3290] = ~(layer_0[10367] ^ layer_0[10593]); 
    assign out[3291] = ~(layer_0[9247] ^ layer_0[9435]); 
    assign out[3292] = layer_0[8142] ^ layer_0[2365]; 
    assign out[3293] = ~(layer_0[6758] ^ layer_0[8742]); 
    assign out[3294] = layer_0[8417] & layer_0[9843]; 
    assign out[3295] = ~(layer_0[10054] | layer_0[11650]); 
    assign out[3296] = ~(layer_0[6626] ^ layer_0[11223]); 
    assign out[3297] = layer_0[5757]; 
    assign out[3298] = layer_0[10806]; 
    assign out[3299] = layer_0[964] ^ layer_0[10971]; 
    assign out[3300] = ~(layer_0[8988] ^ layer_0[2477]); 
    assign out[3301] = ~(layer_0[2018] ^ layer_0[2807]); 
    assign out[3302] = ~(layer_0[1856] ^ layer_0[5438]); 
    assign out[3303] = layer_0[8061]; 
    assign out[3304] = ~layer_0[1825] | (layer_0[1825] & layer_0[887]); 
    assign out[3305] = layer_0[11735] ^ layer_0[8218]; 
    assign out[3306] = layer_0[11783] ^ layer_0[10829]; 
    assign out[3307] = layer_0[1692] ^ layer_0[3281]; 
    assign out[3308] = ~(layer_0[677] ^ layer_0[5650]); 
    assign out[3309] = layer_0[4927] & ~layer_0[4309]; 
    assign out[3310] = layer_0[2983] ^ layer_0[11920]; 
    assign out[3311] = layer_0[1985] ^ layer_0[45]; 
    assign out[3312] = layer_0[947] ^ layer_0[8217]; 
    assign out[3313] = ~(layer_0[2068] & layer_0[7562]); 
    assign out[3314] = layer_0[8391]; 
    assign out[3315] = layer_0[3847] ^ layer_0[4578]; 
    assign out[3316] = ~(layer_0[4317] ^ layer_0[9165]); 
    assign out[3317] = ~layer_0[11184]; 
    assign out[3318] = ~layer_0[9485]; 
    assign out[3319] = ~layer_0[3389]; 
    assign out[3320] = ~layer_0[4941] | (layer_0[4941] & layer_0[10685]); 
    assign out[3321] = layer_0[10115]; 
    assign out[3322] = layer_0[3269] ^ layer_0[8125]; 
    assign out[3323] = ~(layer_0[805] | layer_0[3869]); 
    assign out[3324] = layer_0[3186] | layer_0[2885]; 
    assign out[3325] = ~layer_0[9351]; 
    assign out[3326] = layer_0[5785]; 
    assign out[3327] = layer_0[9415]; 
    assign out[3328] = layer_0[7318] & ~layer_0[647]; 
    assign out[3329] = layer_0[7910] & ~layer_0[11872]; 
    assign out[3330] = layer_0[3336] & ~layer_0[3689]; 
    assign out[3331] = layer_0[4689] & layer_0[6753]; 
    assign out[3332] = ~(layer_0[6319] ^ layer_0[338]); 
    assign out[3333] = ~layer_0[9050]; 
    assign out[3334] = layer_0[10008]; 
    assign out[3335] = layer_0[8058] | layer_0[611]; 
    assign out[3336] = layer_0[1768] ^ layer_0[8722]; 
    assign out[3337] = ~layer_0[10676]; 
    assign out[3338] = ~layer_0[9478]; 
    assign out[3339] = ~(layer_0[10443] ^ layer_0[11984]); 
    assign out[3340] = ~layer_0[3310]; 
    assign out[3341] = layer_0[6398] ^ layer_0[6554]; 
    assign out[3342] = ~layer_0[9184]; 
    assign out[3343] = layer_0[4032] & ~layer_0[2435]; 
    assign out[3344] = layer_0[1715]; 
    assign out[3345] = layer_0[11182] & layer_0[9546]; 
    assign out[3346] = ~(layer_0[10412] ^ layer_0[11220]); 
    assign out[3347] = layer_0[11896] & ~layer_0[11848]; 
    assign out[3348] = layer_0[5682]; 
    assign out[3349] = ~layer_0[69] | (layer_0[69] & layer_0[8149]); 
    assign out[3350] = layer_0[7669]; 
    assign out[3351] = ~(layer_0[11105] ^ layer_0[9031]); 
    assign out[3352] = ~(layer_0[4232] | layer_0[8850]); 
    assign out[3353] = ~(layer_0[1788] ^ layer_0[7627]); 
    assign out[3354] = ~layer_0[4377]; 
    assign out[3355] = ~layer_0[2644]; 
    assign out[3356] = ~(layer_0[1501] ^ layer_0[2059]); 
    assign out[3357] = layer_0[512] ^ layer_0[8767]; 
    assign out[3358] = ~(layer_0[8483] | layer_0[6872]); 
    assign out[3359] = ~layer_0[11312] | (layer_0[11312] & layer_0[6385]); 
    assign out[3360] = ~layer_0[1537]; 
    assign out[3361] = ~(layer_0[9845] ^ layer_0[4860]); 
    assign out[3362] = layer_0[11119] ^ layer_0[3595]; 
    assign out[3363] = layer_0[9131] ^ layer_0[8811]; 
    assign out[3364] = layer_0[4581] ^ layer_0[6651]; 
    assign out[3365] = ~layer_0[1331]; 
    assign out[3366] = layer_0[6017] ^ layer_0[1036]; 
    assign out[3367] = layer_0[9274] & ~layer_0[4671]; 
    assign out[3368] = ~layer_0[5997] | (layer_0[5997] & layer_0[7186]); 
    assign out[3369] = layer_0[1488] ^ layer_0[11795]; 
    assign out[3370] = layer_0[8293]; 
    assign out[3371] = layer_0[11526]; 
    assign out[3372] = ~(layer_0[8654] ^ layer_0[6217]); 
    assign out[3373] = ~layer_0[3753]; 
    assign out[3374] = ~(layer_0[7397] ^ layer_0[4038]); 
    assign out[3375] = ~(layer_0[10011] ^ layer_0[7662]); 
    assign out[3376] = layer_0[3955] & layer_0[9206]; 
    assign out[3377] = layer_0[6400] ^ layer_0[5668]; 
    assign out[3378] = ~(layer_0[10852] ^ layer_0[2544]); 
    assign out[3379] = ~(layer_0[7480] ^ layer_0[236]); 
    assign out[3380] = layer_0[4561] | layer_0[11659]; 
    assign out[3381] = layer_0[9779] ^ layer_0[9197]; 
    assign out[3382] = ~layer_0[7520] | (layer_0[12] & layer_0[7520]); 
    assign out[3383] = ~(layer_0[1386] | layer_0[5186]); 
    assign out[3384] = layer_0[8624] ^ layer_0[2578]; 
    assign out[3385] = ~layer_0[9944] | (layer_0[9944] & layer_0[6715]); 
    assign out[3386] = layer_0[194] ^ layer_0[2033]; 
    assign out[3387] = layer_0[11930] & layer_0[1710]; 
    assign out[3388] = layer_0[230]; 
    assign out[3389] = ~(layer_0[384] ^ layer_0[8864]); 
    assign out[3390] = ~(layer_0[3912] ^ layer_0[3353]); 
    assign out[3391] = ~layer_0[2341]; 
    assign out[3392] = ~(layer_0[7432] ^ layer_0[9850]); 
    assign out[3393] = ~(layer_0[2916] ^ layer_0[2375]); 
    assign out[3394] = ~layer_0[10202] | (layer_0[3091] & layer_0[10202]); 
    assign out[3395] = ~layer_0[7953]; 
    assign out[3396] = ~layer_0[11210] | (layer_0[11210] & layer_0[11033]); 
    assign out[3397] = ~layer_0[5931]; 
    assign out[3398] = ~(layer_0[6656] | layer_0[7817]); 
    assign out[3399] = layer_0[11083] ^ layer_0[115]; 
    assign out[3400] = ~layer_0[6914] | (layer_0[1074] & layer_0[6914]); 
    assign out[3401] = ~(layer_0[11180] | layer_0[4490]); 
    assign out[3402] = layer_0[3124] & ~layer_0[10347]; 
    assign out[3403] = layer_0[2172] & ~layer_0[9262]; 
    assign out[3404] = layer_0[7664] ^ layer_0[8957]; 
    assign out[3405] = layer_0[998] & ~layer_0[9528]; 
    assign out[3406] = ~(layer_0[4047] ^ layer_0[6321]); 
    assign out[3407] = layer_0[4690] & ~layer_0[6440]; 
    assign out[3408] = ~(layer_0[517] | layer_0[1023]); 
    assign out[3409] = ~layer_0[3647] | (layer_0[3647] & layer_0[5565]); 
    assign out[3410] = layer_0[9272] ^ layer_0[2552]; 
    assign out[3411] = layer_0[477] ^ layer_0[7670]; 
    assign out[3412] = layer_0[10389]; 
    assign out[3413] = ~(layer_0[7378] | layer_0[6913]); 
    assign out[3414] = layer_0[1763] & layer_0[7055]; 
    assign out[3415] = ~layer_0[6416]; 
    assign out[3416] = ~(layer_0[3188] ^ layer_0[11536]); 
    assign out[3417] = ~layer_0[5921] | (layer_0[5921] & layer_0[6892]); 
    assign out[3418] = ~layer_0[454]; 
    assign out[3419] = layer_0[6663] & layer_0[9096]; 
    assign out[3420] = ~(layer_0[6253] ^ layer_0[10875]); 
    assign out[3421] = ~(layer_0[8933] | layer_0[688]); 
    assign out[3422] = layer_0[1855] & ~layer_0[9832]; 
    assign out[3423] = ~(layer_0[3673] ^ layer_0[11262]); 
    assign out[3424] = layer_0[8567] ^ layer_0[9720]; 
    assign out[3425] = ~(layer_0[1361] & layer_0[9347]); 
    assign out[3426] = layer_0[3663] ^ layer_0[6331]; 
    assign out[3427] = ~layer_0[2431]; 
    assign out[3428] = layer_0[1464]; 
    assign out[3429] = layer_0[10897] & ~layer_0[9112]; 
    assign out[3430] = layer_0[3111] ^ layer_0[4765]; 
    assign out[3431] = ~(layer_0[2040] ^ layer_0[5376]); 
    assign out[3432] = ~(layer_0[4706] ^ layer_0[5357]); 
    assign out[3433] = layer_0[7990] ^ layer_0[1855]; 
    assign out[3434] = ~(layer_0[1802] ^ layer_0[3650]); 
    assign out[3435] = ~(layer_0[2622] ^ layer_0[6236]); 
    assign out[3436] = layer_0[4527] ^ layer_0[2080]; 
    assign out[3437] = layer_0[322] ^ layer_0[427]; 
    assign out[3438] = layer_0[244] ^ layer_0[9639]; 
    assign out[3439] = layer_0[6691] | layer_0[926]; 
    assign out[3440] = ~(layer_0[10673] ^ layer_0[1096]); 
    assign out[3441] = layer_0[7884] ^ layer_0[398]; 
    assign out[3442] = ~layer_0[1414]; 
    assign out[3443] = layer_0[4128] ^ layer_0[1351]; 
    assign out[3444] = layer_0[3512]; 
    assign out[3445] = layer_0[8237] ^ layer_0[597]; 
    assign out[3446] = layer_0[1974] & ~layer_0[4440]; 
    assign out[3447] = layer_0[1008]; 
    assign out[3448] = layer_0[3581] ^ layer_0[582]; 
    assign out[3449] = ~(layer_0[6386] & layer_0[10483]); 
    assign out[3450] = ~(layer_0[6397] | layer_0[3777]); 
    assign out[3451] = layer_0[7398] & ~layer_0[5297]; 
    assign out[3452] = ~(layer_0[1656] ^ layer_0[10867]); 
    assign out[3453] = ~(layer_0[9640] ^ layer_0[9016]); 
    assign out[3454] = ~(layer_0[8351] ^ layer_0[1353]); 
    assign out[3455] = ~(layer_0[935] ^ layer_0[4669]); 
    assign out[3456] = layer_0[4984]; 
    assign out[3457] = ~(layer_0[6822] | layer_0[6359]); 
    assign out[3458] = ~(layer_0[7233] | layer_0[11134]); 
    assign out[3459] = ~(layer_0[6510] ^ layer_0[10467]); 
    assign out[3460] = layer_0[2700] & ~layer_0[1474]; 
    assign out[3461] = layer_0[8323] ^ layer_0[9807]; 
    assign out[3462] = ~(layer_0[7001] ^ layer_0[7470]); 
    assign out[3463] = ~(layer_0[11357] ^ layer_0[8036]); 
    assign out[3464] = ~(layer_0[4776] ^ layer_0[6824]); 
    assign out[3465] = layer_0[1906]; 
    assign out[3466] = ~(layer_0[8890] ^ layer_0[8776]); 
    assign out[3467] = ~(layer_0[8107] | layer_0[8090]); 
    assign out[3468] = ~layer_0[4097]; 
    assign out[3469] = layer_0[3627] & layer_0[2447]; 
    assign out[3470] = layer_0[6053]; 
    assign out[3471] = ~(layer_0[3211] ^ layer_0[10156]); 
    assign out[3472] = layer_0[11027] ^ layer_0[10473]; 
    assign out[3473] = ~(layer_0[11239] | layer_0[7347]); 
    assign out[3474] = layer_0[611]; 
    assign out[3475] = ~layer_0[3766] | (layer_0[3766] & layer_0[6748]); 
    assign out[3476] = layer_0[6880] ^ layer_0[6388]; 
    assign out[3477] = ~(layer_0[7948] ^ layer_0[5525]); 
    assign out[3478] = layer_0[11808] & layer_0[10377]; 
    assign out[3479] = ~(layer_0[3523] ^ layer_0[4]); 
    assign out[3480] = ~layer_0[8972]; 
    assign out[3481] = layer_0[11380] ^ layer_0[135]; 
    assign out[3482] = ~layer_0[379]; 
    assign out[3483] = layer_0[3657] & ~layer_0[3365]; 
    assign out[3484] = layer_0[9156] ^ layer_0[103]; 
    assign out[3485] = ~(layer_0[2799] ^ layer_0[8623]); 
    assign out[3486] = layer_0[8333] ^ layer_0[5815]; 
    assign out[3487] = ~(layer_0[7125] ^ layer_0[4385]); 
    assign out[3488] = layer_0[10674] ^ layer_0[841]; 
    assign out[3489] = ~(layer_0[2510] ^ layer_0[9636]); 
    assign out[3490] = layer_0[8061] & ~layer_0[4347]; 
    assign out[3491] = layer_0[10522] ^ layer_0[264]; 
    assign out[3492] = ~layer_0[8939]; 
    assign out[3493] = ~layer_0[5605]; 
    assign out[3494] = ~layer_0[6195]; 
    assign out[3495] = ~(layer_0[869] ^ layer_0[6952]); 
    assign out[3496] = layer_0[8497]; 
    assign out[3497] = layer_0[1783]; 
    assign out[3498] = layer_0[11823]; 
    assign out[3499] = layer_0[1874] ^ layer_0[7532]; 
    assign out[3500] = ~(layer_0[2443] ^ layer_0[3683]); 
    assign out[3501] = ~layer_0[1452]; 
    assign out[3502] = layer_0[5117] ^ layer_0[4516]; 
    assign out[3503] = ~(layer_0[5127] ^ layer_0[1357]); 
    assign out[3504] = ~(layer_0[4015] ^ layer_0[3339]); 
    assign out[3505] = ~layer_0[1171] | (layer_0[5857] & layer_0[1171]); 
    assign out[3506] = ~(layer_0[7853] ^ layer_0[10727]); 
    assign out[3507] = layer_0[5405]; 
    assign out[3508] = ~(layer_0[7234] ^ layer_0[7129]); 
    assign out[3509] = ~layer_0[152] | (layer_0[751] & layer_0[152]); 
    assign out[3510] = layer_0[11401] ^ layer_0[1386]; 
    assign out[3511] = layer_0[9738] ^ layer_0[10907]; 
    assign out[3512] = ~layer_0[8034]; 
    assign out[3513] = layer_0[9392] ^ layer_0[4214]; 
    assign out[3514] = ~layer_0[3707]; 
    assign out[3515] = layer_0[4647] ^ layer_0[8770]; 
    assign out[3516] = layer_0[10180] ^ layer_0[8909]; 
    assign out[3517] = ~(layer_0[5654] ^ layer_0[2000]); 
    assign out[3518] = layer_0[8033] & layer_0[3459]; 
    assign out[3519] = ~(layer_0[5741] ^ layer_0[2340]); 
    assign out[3520] = ~layer_0[768]; 
    assign out[3521] = ~(layer_0[2942] ^ layer_0[6803]); 
    assign out[3522] = layer_0[2785] ^ layer_0[11566]; 
    assign out[3523] = layer_0[4356] ^ layer_0[10164]; 
    assign out[3524] = ~layer_0[5614] | (layer_0[5614] & layer_0[9071]); 
    assign out[3525] = layer_0[2845] ^ layer_0[3762]; 
    assign out[3526] = layer_0[9130] & ~layer_0[10832]; 
    assign out[3527] = ~layer_0[8787]; 
    assign out[3528] = ~(layer_0[2338] ^ layer_0[5233]); 
    assign out[3529] = ~(layer_0[11279] ^ layer_0[9232]); 
    assign out[3530] = ~(layer_0[3432] | layer_0[4814]); 
    assign out[3531] = layer_0[3673] & ~layer_0[11391]; 
    assign out[3532] = layer_0[3062]; 
    assign out[3533] = layer_0[3736]; 
    assign out[3534] = layer_0[11133] & layer_0[9355]; 
    assign out[3535] = ~(layer_0[7430] ^ layer_0[1046]); 
    assign out[3536] = layer_0[8004] ^ layer_0[811]; 
    assign out[3537] = layer_0[6098] ^ layer_0[11243]; 
    assign out[3538] = layer_0[8919] & ~layer_0[3210]; 
    assign out[3539] = ~(layer_0[5901] ^ layer_0[3248]); 
    assign out[3540] = ~layer_0[2579]; 
    assign out[3541] = ~(layer_0[6496] ^ layer_0[8791]); 
    assign out[3542] = layer_0[5988] ^ layer_0[3146]; 
    assign out[3543] = ~(layer_0[5651] ^ layer_0[9406]); 
    assign out[3544] = layer_0[1296] ^ layer_0[1167]; 
    assign out[3545] = ~(layer_0[2677] | layer_0[5960]); 
    assign out[3546] = ~(layer_0[10625] ^ layer_0[2398]); 
    assign out[3547] = layer_0[2056] & ~layer_0[5498]; 
    assign out[3548] = layer_0[4705]; 
    assign out[3549] = ~(layer_0[9305] ^ layer_0[8232]); 
    assign out[3550] = ~layer_0[4525]; 
    assign out[3551] = layer_0[5637] & layer_0[2037]; 
    assign out[3552] = ~(layer_0[10162] ^ layer_0[2084]); 
    assign out[3553] = layer_0[9284] & layer_0[2093]; 
    assign out[3554] = layer_0[4962] & ~layer_0[9458]; 
    assign out[3555] = ~layer_0[8257]; 
    assign out[3556] = layer_0[8143] ^ layer_0[10018]; 
    assign out[3557] = layer_0[11337] ^ layer_0[2668]; 
    assign out[3558] = ~layer_0[9431] | (layer_0[2966] & layer_0[9431]); 
    assign out[3559] = layer_0[9679] ^ layer_0[1287]; 
    assign out[3560] = layer_0[658] & layer_0[8575]; 
    assign out[3561] = layer_0[9973]; 
    assign out[3562] = ~(layer_0[9571] ^ layer_0[4045]); 
    assign out[3563] = layer_0[7433] & ~layer_0[2161]; 
    assign out[3564] = ~layer_0[11276]; 
    assign out[3565] = layer_0[2070]; 
    assign out[3566] = layer_0[10475] ^ layer_0[4421]; 
    assign out[3567] = ~(layer_0[2065] | layer_0[11186]); 
    assign out[3568] = layer_0[7880]; 
    assign out[3569] = layer_0[5752] ^ layer_0[7711]; 
    assign out[3570] = ~layer_0[2386] | (layer_0[2386] & layer_0[7220]); 
    assign out[3571] = layer_0[3517] | layer_0[5968]; 
    assign out[3572] = layer_0[3956] | layer_0[11468]; 
    assign out[3573] = ~(layer_0[9391] ^ layer_0[9753]); 
    assign out[3574] = layer_0[2197] | layer_0[9072]; 
    assign out[3575] = layer_0[5972]; 
    assign out[3576] = ~(layer_0[721] ^ layer_0[2604]); 
    assign out[3577] = ~(layer_0[8240] | layer_0[10210]); 
    assign out[3578] = layer_0[7298]; 
    assign out[3579] = ~layer_0[3164]; 
    assign out[3580] = layer_0[11202] & ~layer_0[2736]; 
    assign out[3581] = layer_0[1163] & ~layer_0[11130]; 
    assign out[3582] = layer_0[663] ^ layer_0[6073]; 
    assign out[3583] = ~layer_0[2587]; 
    assign out[3584] = layer_0[11001] ^ layer_0[1452]; 
    assign out[3585] = ~(layer_0[4365] ^ layer_0[9489]); 
    assign out[3586] = ~(layer_0[6039] ^ layer_0[1506]); 
    assign out[3587] = layer_0[2803] ^ layer_0[7317]; 
    assign out[3588] = ~layer_0[7885]; 
    assign out[3589] = layer_0[9522] ^ layer_0[1918]; 
    assign out[3590] = layer_0[8262] ^ layer_0[5821]; 
    assign out[3591] = ~(layer_0[6192] ^ layer_0[3450]); 
    assign out[3592] = ~(layer_0[11145] ^ layer_0[9883]); 
    assign out[3593] = ~(layer_0[2656] | layer_0[746]); 
    assign out[3594] = layer_0[9374] ^ layer_0[5588]; 
    assign out[3595] = ~(layer_0[11992] | layer_0[3903]); 
    assign out[3596] = layer_0[1398] ^ layer_0[11419]; 
    assign out[3597] = layer_0[11569] ^ layer_0[4626]; 
    assign out[3598] = ~(layer_0[8744] | layer_0[7286]); 
    assign out[3599] = ~(layer_0[8239] ^ layer_0[156]); 
    assign out[3600] = layer_0[5977] ^ layer_0[10177]; 
    assign out[3601] = ~(layer_0[223] | layer_0[9105]); 
    assign out[3602] = ~layer_0[5276]; 
    assign out[3603] = ~layer_0[9981] | (layer_0[11551] & layer_0[9981]); 
    assign out[3604] = layer_0[1062] ^ layer_0[11879]; 
    assign out[3605] = layer_0[886] ^ layer_0[8765]; 
    assign out[3606] = ~(layer_0[7781] ^ layer_0[3098]); 
    assign out[3607] = ~layer_0[2065]; 
    assign out[3608] = layer_0[6277] & ~layer_0[9794]; 
    assign out[3609] = ~(layer_0[7431] ^ layer_0[7565]); 
    assign out[3610] = ~(layer_0[11705] ^ layer_0[4104]); 
    assign out[3611] = layer_0[2468] & ~layer_0[1622]; 
    assign out[3612] = layer_0[6084] ^ layer_0[243]; 
    assign out[3613] = layer_0[3727]; 
    assign out[3614] = ~(layer_0[1138] ^ layer_0[3845]); 
    assign out[3615] = ~(layer_0[999] | layer_0[11418]); 
    assign out[3616] = layer_0[8218] ^ layer_0[9614]; 
    assign out[3617] = ~(layer_0[5439] ^ layer_0[9147]); 
    assign out[3618] = layer_0[5928] ^ layer_0[6114]; 
    assign out[3619] = ~(layer_0[879] & layer_0[884]); 
    assign out[3620] = layer_0[1689]; 
    assign out[3621] = layer_0[7094]; 
    assign out[3622] = ~(layer_0[3150] | layer_0[9331]); 
    assign out[3623] = layer_0[6235]; 
    assign out[3624] = layer_0[11654] ^ layer_0[9462]; 
    assign out[3625] = ~layer_0[11658]; 
    assign out[3626] = ~(layer_0[2003] ^ layer_0[4408]); 
    assign out[3627] = ~(layer_0[9724] ^ layer_0[9877]); 
    assign out[3628] = ~layer_0[7934] | (layer_0[7934] & layer_0[6493]); 
    assign out[3629] = ~(layer_0[9162] ^ layer_0[7007]); 
    assign out[3630] = ~layer_0[9121]; 
    assign out[3631] = layer_0[2428] ^ layer_0[5927]; 
    assign out[3632] = ~layer_0[7603]; 
    assign out[3633] = ~(layer_0[8120] ^ layer_0[5067]); 
    assign out[3634] = ~layer_0[2146]; 
    assign out[3635] = layer_0[6522] | layer_0[6640]; 
    assign out[3636] = layer_0[9900] ^ layer_0[2727]; 
    assign out[3637] = ~layer_0[5373] | (layer_0[5373] & layer_0[6285]); 
    assign out[3638] = ~(layer_0[11493] ^ layer_0[4246]); 
    assign out[3639] = ~(layer_0[9809] ^ layer_0[11288]); 
    assign out[3640] = layer_0[4940] ^ layer_0[10286]; 
    assign out[3641] = layer_0[3953] & ~layer_0[5430]; 
    assign out[3642] = layer_0[8469] ^ layer_0[1813]; 
    assign out[3643] = ~(layer_0[11442] ^ layer_0[10614]); 
    assign out[3644] = layer_0[2] ^ layer_0[4294]; 
    assign out[3645] = layer_0[4604] & ~layer_0[10634]; 
    assign out[3646] = ~(layer_0[2553] | layer_0[3487]); 
    assign out[3647] = layer_0[3121] ^ layer_0[3931]; 
    assign out[3648] = layer_0[10641] ^ layer_0[4719]; 
    assign out[3649] = ~(layer_0[7126] ^ layer_0[9211]); 
    assign out[3650] = layer_0[4341] ^ layer_0[3021]; 
    assign out[3651] = layer_0[1218] & ~layer_0[5502]; 
    assign out[3652] = layer_0[8550] ^ layer_0[5128]; 
    assign out[3653] = ~(layer_0[10439] ^ layer_0[9893]); 
    assign out[3654] = ~(layer_0[9604] ^ layer_0[7185]); 
    assign out[3655] = ~(layer_0[10579] ^ layer_0[263]); 
    assign out[3656] = layer_0[11692] ^ layer_0[5045]; 
    assign out[3657] = ~(layer_0[1643] ^ layer_0[11381]); 
    assign out[3658] = ~(layer_0[9321] ^ layer_0[7419]); 
    assign out[3659] = ~(layer_0[3851] | layer_0[8236]); 
    assign out[3660] = ~(layer_0[11496] ^ layer_0[7791]); 
    assign out[3661] = layer_0[4475] ^ layer_0[5699]; 
    assign out[3662] = layer_0[2640] & ~layer_0[3332]; 
    assign out[3663] = layer_0[6361]; 
    assign out[3664] = ~(layer_0[6137] | layer_0[2060]); 
    assign out[3665] = ~layer_0[1553] | (layer_0[1553] & layer_0[3546]); 
    assign out[3666] = layer_0[7547] & ~layer_0[6889]; 
    assign out[3667] = layer_0[3257] & layer_0[10394]; 
    assign out[3668] = layer_0[1747] & ~layer_0[8013]; 
    assign out[3669] = layer_0[11385] & ~layer_0[6723]; 
    assign out[3670] = ~layer_0[10630]; 
    assign out[3671] = ~(layer_0[6357] ^ layer_0[7095]); 
    assign out[3672] = layer_0[6567]; 
    assign out[3673] = layer_0[2775] | layer_0[7541]; 
    assign out[3674] = layer_0[11994]; 
    assign out[3675] = ~layer_0[11633]; 
    assign out[3676] = layer_0[7668] ^ layer_0[6995]; 
    assign out[3677] = ~(layer_0[9475] | layer_0[122]); 
    assign out[3678] = layer_0[9330] ^ layer_0[9187]; 
    assign out[3679] = ~(layer_0[389] ^ layer_0[10894]); 
    assign out[3680] = ~(layer_0[2165] ^ layer_0[10905]); 
    assign out[3681] = layer_0[7145]; 
    assign out[3682] = layer_0[447] ^ layer_0[1636]; 
    assign out[3683] = layer_0[8479] ^ layer_0[9189]; 
    assign out[3684] = layer_0[2618] & ~layer_0[1364]; 
    assign out[3685] = ~(layer_0[77] ^ layer_0[11857]); 
    assign out[3686] = layer_0[3323] ^ layer_0[10776]; 
    assign out[3687] = layer_0[10870] & ~layer_0[1471]; 
    assign out[3688] = ~layer_0[2498] | (layer_0[9659] & layer_0[2498]); 
    assign out[3689] = ~(layer_0[6402] ^ layer_0[8671]); 
    assign out[3690] = layer_0[10444] ^ layer_0[6326]; 
    assign out[3691] = ~(layer_0[6797] | layer_0[4830]); 
    assign out[3692] = layer_0[4165] ^ layer_0[4402]; 
    assign out[3693] = layer_0[4035] ^ layer_0[4194]; 
    assign out[3694] = ~(layer_0[9903] | layer_0[5783]); 
    assign out[3695] = ~(layer_0[1055] ^ layer_0[1623]); 
    assign out[3696] = ~(layer_0[9303] & layer_0[385]); 
    assign out[3697] = layer_0[7586] & ~layer_0[1544]; 
    assign out[3698] = layer_0[10071] & ~layer_0[2722]; 
    assign out[3699] = ~(layer_0[5130] ^ layer_0[7422]); 
    assign out[3700] = layer_0[2799] ^ layer_0[7218]; 
    assign out[3701] = layer_0[593] ^ layer_0[11763]; 
    assign out[3702] = ~layer_0[9965]; 
    assign out[3703] = layer_0[1209] ^ layer_0[11598]; 
    assign out[3704] = ~(layer_0[4085] ^ layer_0[11193]); 
    assign out[3705] = ~(layer_0[3065] ^ layer_0[10306]); 
    assign out[3706] = layer_0[1783] ^ layer_0[6875]; 
    assign out[3707] = layer_0[2600]; 
    assign out[3708] = ~(layer_0[10758] ^ layer_0[11955]); 
    assign out[3709] = ~layer_0[3155]; 
    assign out[3710] = layer_0[5090]; 
    assign out[3711] = layer_0[10445] ^ layer_0[4513]; 
    assign out[3712] = ~(layer_0[3014] | layer_0[4279]); 
    assign out[3713] = layer_0[5050] & ~layer_0[8941]; 
    assign out[3714] = ~(layer_0[1174] ^ layer_0[11773]); 
    assign out[3715] = layer_0[4815] ^ layer_0[10964]; 
    assign out[3716] = layer_0[10181] ^ layer_0[361]; 
    assign out[3717] = ~(layer_0[8141] ^ layer_0[6169]); 
    assign out[3718] = ~layer_0[5711]; 
    assign out[3719] = layer_0[7240] & ~layer_0[7197]; 
    assign out[3720] = layer_0[2735] ^ layer_0[7618]; 
    assign out[3721] = layer_0[3736] & layer_0[129]; 
    assign out[3722] = ~layer_0[8478]; 
    assign out[3723] = layer_0[7746]; 
    assign out[3724] = ~(layer_0[6236] ^ layer_0[8872]); 
    assign out[3725] = ~(layer_0[10062] ^ layer_0[2633]); 
    assign out[3726] = ~(layer_0[2238] | layer_0[11484]); 
    assign out[3727] = layer_0[6637] ^ layer_0[2137]; 
    assign out[3728] = ~(layer_0[1620] ^ layer_0[1034]); 
    assign out[3729] = ~(layer_0[10203] | layer_0[9794]); 
    assign out[3730] = ~layer_0[7030]; 
    assign out[3731] = layer_0[1905] & ~layer_0[5331]; 
    assign out[3732] = ~(layer_0[279] ^ layer_0[7426]); 
    assign out[3733] = layer_0[4213]; 
    assign out[3734] = ~(layer_0[1415] & layer_0[5460]); 
    assign out[3735] = layer_0[6986] ^ layer_0[4681]; 
    assign out[3736] = layer_0[472]; 
    assign out[3737] = ~(layer_0[8690] ^ layer_0[4715]); 
    assign out[3738] = ~layer_0[6551] | (layer_0[10698] & layer_0[6551]); 
    assign out[3739] = ~layer_0[2305] | (layer_0[9524] & layer_0[2305]); 
    assign out[3740] = layer_0[8754] ^ layer_0[2466]; 
    assign out[3741] = layer_0[748]; 
    assign out[3742] = ~(layer_0[9467] ^ layer_0[7457]); 
    assign out[3743] = ~layer_0[7837] | (layer_0[7232] & layer_0[7837]); 
    assign out[3744] = ~(layer_0[441] ^ layer_0[8597]); 
    assign out[3745] = ~(layer_0[10339] ^ layer_0[11084]); 
    assign out[3746] = layer_0[3130]; 
    assign out[3747] = ~(layer_0[7279] ^ layer_0[10370]); 
    assign out[3748] = ~layer_0[9927] | (layer_0[9927] & layer_0[2875]); 
    assign out[3749] = ~(layer_0[4036] ^ layer_0[6343]); 
    assign out[3750] = ~(layer_0[4260] ^ layer_0[5328]); 
    assign out[3751] = layer_0[8807] | layer_0[11826]; 
    assign out[3752] = layer_0[11364] ^ layer_0[5570]; 
    assign out[3753] = ~(layer_0[5643] ^ layer_0[2053]); 
    assign out[3754] = ~(layer_0[3197] & layer_0[2004]); 
    assign out[3755] = layer_0[9655] & ~layer_0[474]; 
    assign out[3756] = layer_0[7769] ^ layer_0[1605]; 
    assign out[3757] = layer_0[4252] ^ layer_0[8156]; 
    assign out[3758] = ~(layer_0[6624] ^ layer_0[9837]); 
    assign out[3759] = ~(layer_0[4886] ^ layer_0[10435]); 
    assign out[3760] = layer_0[681] & ~layer_0[1953]; 
    assign out[3761] = layer_0[2997] & ~layer_0[1331]; 
    assign out[3762] = layer_0[91]; 
    assign out[3763] = layer_0[1526] & layer_0[4366]; 
    assign out[3764] = layer_0[3825]; 
    assign out[3765] = layer_0[5353] & ~layer_0[4333]; 
    assign out[3766] = layer_0[11232] ^ layer_0[4446]; 
    assign out[3767] = layer_0[5716] ^ layer_0[11496]; 
    assign out[3768] = ~(layer_0[11393] ^ layer_0[7395]); 
    assign out[3769] = layer_0[6119] ^ layer_0[7987]; 
    assign out[3770] = layer_0[7307] ^ layer_0[4164]; 
    assign out[3771] = ~(layer_0[4763] ^ layer_0[7833]); 
    assign out[3772] = ~(layer_0[1075] & layer_0[1402]); 
    assign out[3773] = layer_0[8609] ^ layer_0[9614]; 
    assign out[3774] = ~(layer_0[10694] | layer_0[8813]); 
    assign out[3775] = ~(layer_0[3158] ^ layer_0[7726]); 
    assign out[3776] = ~(layer_0[11906] ^ layer_0[5112]); 
    assign out[3777] = ~(layer_0[1010] | layer_0[6291]); 
    assign out[3778] = ~(layer_0[7868] ^ layer_0[3894]); 
    assign out[3779] = layer_0[5953] ^ layer_0[4778]; 
    assign out[3780] = ~(layer_0[11444] ^ layer_0[453]); 
    assign out[3781] = ~(layer_0[862] ^ layer_0[6908]); 
    assign out[3782] = layer_0[2836] ^ layer_0[9534]; 
    assign out[3783] = layer_0[6851]; 
    assign out[3784] = layer_0[4722]; 
    assign out[3785] = ~layer_0[1691]; 
    assign out[3786] = ~(layer_0[9196] ^ layer_0[1066]); 
    assign out[3787] = layer_0[3856] & layer_0[5162]; 
    assign out[3788] = ~(layer_0[4316] ^ layer_0[4494]); 
    assign out[3789] = layer_0[4221]; 
    assign out[3790] = layer_0[5337] & layer_0[1777]; 
    assign out[3791] = layer_0[1307]; 
    assign out[3792] = ~(layer_0[838] ^ layer_0[5624]); 
    assign out[3793] = ~layer_0[383]; 
    assign out[3794] = ~(layer_0[4302] | layer_0[6382]); 
    assign out[3795] = layer_0[7365]; 
    assign out[3796] = ~(layer_0[3884] ^ layer_0[7749]); 
    assign out[3797] = ~layer_0[4863]; 
    assign out[3798] = ~layer_0[1009]; 
    assign out[3799] = layer_0[6098]; 
    assign out[3800] = ~(layer_0[3172] ^ layer_0[6525]); 
    assign out[3801] = ~layer_0[9654]; 
    assign out[3802] = layer_0[7066] & ~layer_0[2333]; 
    assign out[3803] = layer_0[4335] ^ layer_0[6132]; 
    assign out[3804] = layer_0[3518] ^ layer_0[8093]; 
    assign out[3805] = layer_0[1128]; 
    assign out[3806] = ~(layer_0[8403] ^ layer_0[2449]); 
    assign out[3807] = ~(layer_0[11407] ^ layer_0[6108]); 
    assign out[3808] = ~layer_0[9906]; 
    assign out[3809] = layer_0[10081] & ~layer_0[340]; 
    assign out[3810] = layer_0[3688]; 
    assign out[3811] = layer_0[7410] & ~layer_0[9813]; 
    assign out[3812] = layer_0[8752] ^ layer_0[316]; 
    assign out[3813] = ~layer_0[577]; 
    assign out[3814] = layer_0[9498] ^ layer_0[5652]; 
    assign out[3815] = layer_0[11497] & ~layer_0[8769]; 
    assign out[3816] = layer_0[7741] ^ layer_0[6387]; 
    assign out[3817] = ~(layer_0[5303] | layer_0[754]); 
    assign out[3818] = layer_0[7870] ^ layer_0[3831]; 
    assign out[3819] = ~layer_0[2756]; 
    assign out[3820] = layer_0[8839]; 
    assign out[3821] = layer_0[5053] ^ layer_0[10800]; 
    assign out[3822] = layer_0[5440] ^ layer_0[5366]; 
    assign out[3823] = ~(layer_0[11899] ^ layer_0[2359]); 
    assign out[3824] = layer_0[9052] & ~layer_0[6617]; 
    assign out[3825] = layer_0[7040] & ~layer_0[3272]; 
    assign out[3826] = layer_0[1245]; 
    assign out[3827] = layer_0[642] ^ layer_0[7031]; 
    assign out[3828] = layer_0[8124]; 
    assign out[3829] = layer_0[6606] & ~layer_0[6568]; 
    assign out[3830] = ~(layer_0[763] ^ layer_0[1815]); 
    assign out[3831] = ~(layer_0[6794] | layer_0[4369]); 
    assign out[3832] = layer_0[943]; 
    assign out[3833] = layer_0[6045] & layer_0[1333]; 
    assign out[3834] = ~(layer_0[6912] & layer_0[11007]); 
    assign out[3835] = layer_0[8187] ^ layer_0[10145]; 
    assign out[3836] = layer_0[9631] & ~layer_0[7605]; 
    assign out[3837] = ~(layer_0[7731] | layer_0[1298]); 
    assign out[3838] = ~layer_0[4134]; 
    assign out[3839] = ~(layer_0[9357] ^ layer_0[8078]); 
    assign out[3840] = ~layer_0[9783] | (layer_0[1646] & layer_0[9783]); 
    assign out[3841] = layer_0[5660]; 
    assign out[3842] = layer_0[6212] & layer_0[3380]; 
    assign out[3843] = ~(layer_0[2821] ^ layer_0[2906]); 
    assign out[3844] = layer_0[9269]; 
    assign out[3845] = ~(layer_0[5945] ^ layer_0[548]); 
    assign out[3846] = ~(layer_0[6699] ^ layer_0[11302]); 
    assign out[3847] = layer_0[10190] ^ layer_0[9078]; 
    assign out[3848] = layer_0[3418] ^ layer_0[6975]; 
    assign out[3849] = layer_0[3774] ^ layer_0[1510]; 
    assign out[3850] = layer_0[8314] ^ layer_0[5805]; 
    assign out[3851] = ~(layer_0[6634] ^ layer_0[9414]); 
    assign out[3852] = layer_0[6595]; 
    assign out[3853] = ~(layer_0[514] ^ layer_0[9750]); 
    assign out[3854] = ~layer_0[7128]; 
    assign out[3855] = layer_0[9289]; 
    assign out[3856] = layer_0[3650] & layer_0[7179]; 
    assign out[3857] = ~(layer_0[10141] & layer_0[1771]); 
    assign out[3858] = layer_0[8402] ^ layer_0[10103]; 
    assign out[3859] = layer_0[9452]; 
    assign out[3860] = layer_0[338] ^ layer_0[9517]; 
    assign out[3861] = ~(layer_0[6870] ^ layer_0[9295]); 
    assign out[3862] = layer_0[1726]; 
    assign out[3863] = layer_0[9279] ^ layer_0[739]; 
    assign out[3864] = layer_0[11103] ^ layer_0[1645]; 
    assign out[3865] = layer_0[4756] & ~layer_0[5483]; 
    assign out[3866] = ~(layer_0[950] ^ layer_0[7263]); 
    assign out[3867] = layer_0[7679] & ~layer_0[10564]; 
    assign out[3868] = ~(layer_0[8833] ^ layer_0[4593]); 
    assign out[3869] = layer_0[4040] & ~layer_0[11363]; 
    assign out[3870] = ~(layer_0[8870] ^ layer_0[10756]); 
    assign out[3871] = layer_0[4705]; 
    assign out[3872] = layer_0[5996]; 
    assign out[3873] = ~(layer_0[8880] ^ layer_0[2421]); 
    assign out[3874] = layer_0[7491] & ~layer_0[9921]; 
    assign out[3875] = layer_0[1254] & layer_0[5584]; 
    assign out[3876] = ~(layer_0[1813] ^ layer_0[7246]); 
    assign out[3877] = ~(layer_0[5245] ^ layer_0[11060]); 
    assign out[3878] = ~(layer_0[7026] ^ layer_0[3358]); 
    assign out[3879] = ~(layer_0[2033] ^ layer_0[2826]); 
    assign out[3880] = ~(layer_0[6694] ^ layer_0[1460]); 
    assign out[3881] = layer_0[6128] ^ layer_0[6651]; 
    assign out[3882] = ~(layer_0[8681] ^ layer_0[999]); 
    assign out[3883] = ~(layer_0[1175] ^ layer_0[2898]); 
    assign out[3884] = layer_0[1652] ^ layer_0[1883]; 
    assign out[3885] = ~(layer_0[538] ^ layer_0[422]); 
    assign out[3886] = ~(layer_0[8904] ^ layer_0[6210]); 
    assign out[3887] = ~layer_0[3103]; 
    assign out[3888] = ~(layer_0[10843] ^ layer_0[11844]); 
    assign out[3889] = ~(layer_0[5683] ^ layer_0[6665]); 
    assign out[3890] = layer_0[7780] ^ layer_0[2307]; 
    assign out[3891] = ~(layer_0[8067] ^ layer_0[175]); 
    assign out[3892] = ~(layer_0[6254] ^ layer_0[784]); 
    assign out[3893] = ~(layer_0[11523] ^ layer_0[10299]); 
    assign out[3894] = layer_0[11090]; 
    assign out[3895] = layer_0[3793]; 
    assign out[3896] = ~layer_0[2521]; 
    assign out[3897] = layer_0[5531] & ~layer_0[4027]; 
    assign out[3898] = ~(layer_0[554] ^ layer_0[6850]); 
    assign out[3899] = ~(layer_0[1037] ^ layer_0[8777]); 
    assign out[3900] = layer_0[6317]; 
    assign out[3901] = ~(layer_0[246] | layer_0[7829]); 
    assign out[3902] = layer_0[8537] ^ layer_0[5464]; 
    assign out[3903] = layer_0[11909] ^ layer_0[4687]; 
    assign out[3904] = layer_0[4058] & ~layer_0[8412]; 
    assign out[3905] = layer_0[6779] ^ layer_0[6103]; 
    assign out[3906] = ~layer_0[3423] | (layer_0[3423] & layer_0[3214]); 
    assign out[3907] = ~layer_0[188] | (layer_0[188] & layer_0[2231]); 
    assign out[3908] = layer_0[3008] ^ layer_0[4239]; 
    assign out[3909] = layer_0[4963]; 
    assign out[3910] = layer_0[6395] & ~layer_0[11191]; 
    assign out[3911] = ~(layer_0[11517] ^ layer_0[11137]); 
    assign out[3912] = layer_0[7925] & ~layer_0[11108]; 
    assign out[3913] = layer_0[1618] ^ layer_0[10098]; 
    assign out[3914] = layer_0[4472] ^ layer_0[6263]; 
    assign out[3915] = ~layer_0[59]; 
    assign out[3916] = ~(layer_0[8110] | layer_0[10854]); 
    assign out[3917] = ~(layer_0[6478] ^ layer_0[9434]); 
    assign out[3918] = ~(layer_0[11402] ^ layer_0[5168]); 
    assign out[3919] = layer_0[5558] & ~layer_0[2184]; 
    assign out[3920] = ~(layer_0[6630] | layer_0[2053]); 
    assign out[3921] = ~layer_0[8084]; 
    assign out[3922] = ~(layer_0[5943] ^ layer_0[4849]); 
    assign out[3923] = layer_0[9451] | layer_0[8472]; 
    assign out[3924] = ~(layer_0[5057] ^ layer_0[4320]); 
    assign out[3925] = ~layer_0[8473]; 
    assign out[3926] = ~(layer_0[5801] ^ layer_0[2289]); 
    assign out[3927] = ~(layer_0[8338] ^ layer_0[3586]); 
    assign out[3928] = ~(layer_0[2362] ^ layer_0[8277]); 
    assign out[3929] = ~(layer_0[7382] ^ layer_0[6796]); 
    assign out[3930] = layer_0[11101] & layer_0[4329]; 
    assign out[3931] = layer_0[9571] ^ layer_0[226]; 
    assign out[3932] = layer_0[8176]; 
    assign out[3933] = layer_0[2226] & ~layer_0[8358]; 
    assign out[3934] = ~(layer_0[8665] ^ layer_0[5187]); 
    assign out[3935] = ~layer_0[9868]; 
    assign out[3936] = layer_0[3302] ^ layer_0[6476]; 
    assign out[3937] = ~(layer_0[6648] ^ layer_0[10992]); 
    assign out[3938] = layer_0[6128] ^ layer_0[1771]; 
    assign out[3939] = layer_0[10787] ^ layer_0[308]; 
    assign out[3940] = layer_0[6885]; 
    assign out[3941] = layer_0[3196] | layer_0[9818]; 
    assign out[3942] = layer_0[4363] ^ layer_0[147]; 
    assign out[3943] = layer_0[9801] ^ layer_0[6608]; 
    assign out[3944] = layer_0[8528]; 
    assign out[3945] = layer_0[8113] ^ layer_0[831]; 
    assign out[3946] = ~(layer_0[4449] ^ layer_0[2471]); 
    assign out[3947] = layer_0[8823]; 
    assign out[3948] = ~layer_0[7487] | (layer_0[11362] & layer_0[7487]); 
    assign out[3949] = ~(layer_0[6247] ^ layer_0[10213]); 
    assign out[3950] = layer_0[5680] ^ layer_0[3679]; 
    assign out[3951] = ~(layer_0[4642] ^ layer_0[7260]); 
    assign out[3952] = ~(layer_0[6322] ^ layer_0[4906]); 
    assign out[3953] = ~(layer_0[6358] ^ layer_0[2768]); 
    assign out[3954] = layer_0[1750]; 
    assign out[3955] = layer_0[8263] & layer_0[11726]; 
    assign out[3956] = layer_0[693] & layer_0[9680]; 
    assign out[3957] = layer_0[7046] ^ layer_0[1478]; 
    assign out[3958] = layer_0[979] & ~layer_0[7219]; 
    assign out[3959] = layer_0[5692]; 
    assign out[3960] = ~layer_0[7981]; 
    assign out[3961] = layer_0[11530] ^ layer_0[190]; 
    assign out[3962] = layer_0[11843] & ~layer_0[9760]; 
    assign out[3963] = ~(layer_0[10015] ^ layer_0[9697]); 
    assign out[3964] = ~(layer_0[6268] ^ layer_0[9303]); 
    assign out[3965] = layer_0[8171] & ~layer_0[8327]; 
    assign out[3966] = layer_0[10076]; 
    assign out[3967] = layer_0[1958]; 
    assign out[3968] = ~(layer_0[8563] ^ layer_0[11586]); 
    assign out[3969] = ~layer_0[1085]; 
    assign out[3970] = ~(layer_0[3996] ^ layer_0[6449]); 
    assign out[3971] = layer_0[11072] & layer_0[6658]; 
    assign out[3972] = ~(layer_0[5407] ^ layer_0[9869]); 
    assign out[3973] = ~layer_0[8053] | (layer_0[4522] & layer_0[8053]); 
    assign out[3974] = ~(layer_0[5975] ^ layer_0[1234]); 
    assign out[3975] = ~(layer_0[7537] ^ layer_0[11722]); 
    assign out[3976] = ~(layer_0[8302] ^ layer_0[5185]); 
    assign out[3977] = ~(layer_0[551] ^ layer_0[10144]); 
    assign out[3978] = layer_0[8984] ^ layer_0[6381]; 
    assign out[3979] = ~(layer_0[7551] ^ layer_0[2548]); 
    assign out[3980] = ~layer_0[8615]; 
    assign out[3981] = layer_0[9451]; 
    assign out[3982] = ~(layer_0[8676] | layer_0[4355]); 
    assign out[3983] = ~layer_0[11116] | (layer_0[11116] & layer_0[4074]); 
    assign out[3984] = layer_0[2030] ^ layer_0[8916]; 
    assign out[3985] = layer_0[6638] & ~layer_0[7473]; 
    assign out[3986] = ~(layer_0[7427] | layer_0[10193]); 
    assign out[3987] = layer_0[4376] ^ layer_0[2977]; 
    assign out[3988] = layer_0[3816]; 
    assign out[3989] = ~(layer_0[2318] ^ layer_0[6594]); 
    assign out[3990] = ~(layer_0[7242] ^ layer_0[9796]); 
    assign out[3991] = layer_0[8571] ^ layer_0[6038]; 
    assign out[3992] = layer_0[5829] ^ layer_0[9865]; 
    assign out[3993] = layer_0[4151] ^ layer_0[224]; 
    assign out[3994] = layer_0[1574] ^ layer_0[2511]; 
    assign out[3995] = ~layer_0[8893]; 
    assign out[3996] = layer_0[526] ^ layer_0[7501]; 
    assign out[3997] = ~(layer_0[10588] ^ layer_0[8991]); 
    assign out[3998] = layer_0[11022] & ~layer_0[1181]; 
    assign out[3999] = ~(layer_0[5486] | layer_0[4257]); 
    assign out[4000] = layer_0[823] | layer_0[10876]; 
    assign out[4001] = layer_0[4073]; 
    assign out[4002] = layer_0[3320] & ~layer_0[8139]; 
    assign out[4003] = layer_0[5006]; 
    assign out[4004] = layer_0[9265] & ~layer_0[3347]; 
    assign out[4005] = layer_0[9675] & layer_0[4203]; 
    assign out[4006] = ~(layer_0[4322] ^ layer_0[6633]); 
    assign out[4007] = layer_0[10545] ^ layer_0[8549]; 
    assign out[4008] = ~layer_0[7235]; 
    assign out[4009] = ~layer_0[6863]; 
    assign out[4010] = layer_0[1201]; 
    assign out[4011] = ~(layer_0[5606] ^ layer_0[2310]); 
    assign out[4012] = layer_0[7139] | layer_0[6430]; 
    assign out[4013] = layer_0[3934] ^ layer_0[5362]; 
    assign out[4014] = ~(layer_0[10857] ^ layer_0[4754]); 
    assign out[4015] = layer_0[3122] ^ layer_0[10065]; 
    assign out[4016] = ~layer_0[4810] | (layer_0[3964] & layer_0[4810]); 
    assign out[4017] = layer_0[1111] ^ layer_0[3883]; 
    assign out[4018] = ~(layer_0[2082] & layer_0[7782]); 
    assign out[4019] = ~(layer_0[146] | layer_0[9318]); 
    assign out[4020] = ~(layer_0[5910] & layer_0[2253]); 
    assign out[4021] = layer_0[5812] ^ layer_0[10192]; 
    assign out[4022] = layer_0[9908] ^ layer_0[8335]; 
    assign out[4023] = layer_0[5856] & ~layer_0[11318]; 
    assign out[4024] = layer_0[6170] | layer_0[6308]; 
    assign out[4025] = layer_0[8345] & ~layer_0[3965]; 
    assign out[4026] = ~layer_0[10848]; 
    assign out[4027] = ~(layer_0[4103] & layer_0[3957]); 
    assign out[4028] = layer_0[1573]; 
    assign out[4029] = layer_0[876] ^ layer_0[3646]; 
    assign out[4030] = ~layer_0[5919]; 
    assign out[4031] = layer_0[10120]; 
    assign out[4032] = ~layer_0[3465] | (layer_0[3465] & layer_0[1274]); 
    assign out[4033] = ~(layer_0[5164] | layer_0[1915]); 
    assign out[4034] = layer_0[2426]; 
    assign out[4035] = ~(layer_0[649] & layer_0[2584]); 
    assign out[4036] = ~layer_0[10388] | (layer_0[10388] & layer_0[4926]); 
    assign out[4037] = layer_0[1844]; 
    assign out[4038] = ~(layer_0[4195] ^ layer_0[1303]); 
    assign out[4039] = layer_0[6785] ^ layer_0[2528]; 
    assign out[4040] = ~(layer_0[3704] ^ layer_0[10865]); 
    assign out[4041] = ~(layer_0[4443] & layer_0[10956]); 
    assign out[4042] = layer_0[4209] ^ layer_0[5355]; 
    assign out[4043] = layer_0[9225] | layer_0[3680]; 
    assign out[4044] = ~(layer_0[8913] & layer_0[1435]); 
    assign out[4045] = ~layer_0[8705]; 
    assign out[4046] = ~(layer_0[6214] ^ layer_0[9939]); 
    assign out[4047] = layer_0[5790]; 
    assign out[4048] = layer_0[6923]; 
    assign out[4049] = ~(layer_0[9437] ^ layer_0[4893]); 
    assign out[4050] = ~layer_0[4849] | (layer_0[4905] & layer_0[4849]); 
    assign out[4051] = ~layer_0[7372] | (layer_0[7372] & layer_0[8667]); 
    assign out[4052] = layer_0[2998] | layer_0[1070]; 
    assign out[4053] = layer_0[6337] ^ layer_0[4401]; 
    assign out[4054] = ~layer_0[5789]; 
    assign out[4055] = ~layer_0[6557] | (layer_0[2406] & layer_0[6557]); 
    assign out[4056] = layer_0[4710] ^ layer_0[3368]; 
    assign out[4057] = layer_0[435] ^ layer_0[3624]; 
    assign out[4058] = layer_0[2854]; 
    assign out[4059] = layer_0[7226] ^ layer_0[7166]; 
    assign out[4060] = ~layer_0[7891] | (layer_0[7891] & layer_0[8648]); 
    assign out[4061] = layer_0[109] | layer_0[8274]; 
    assign out[4062] = ~(layer_0[2019] ^ layer_0[4628]); 
    assign out[4063] = layer_0[4471] & layer_0[8280]; 
    assign out[4064] = ~(layer_0[1361] & layer_0[3409]); 
    assign out[4065] = ~layer_0[4196] | (layer_0[4861] & layer_0[4196]); 
    assign out[4066] = ~layer_0[7906] | (layer_0[9495] & layer_0[7906]); 
    assign out[4067] = layer_0[6575] ^ layer_0[11273]; 
    assign out[4068] = ~(layer_0[762] ^ layer_0[3592]); 
    assign out[4069] = ~layer_0[8731] | (layer_0[8731] & layer_0[10516]); 
    assign out[4070] = ~layer_0[833]; 
    assign out[4071] = ~layer_0[6091] | (layer_0[6091] & layer_0[3173]); 
    assign out[4072] = layer_0[2487]; 
    assign out[4073] = ~(layer_0[3270] ^ layer_0[6951]); 
    assign out[4074] = ~layer_0[2422] | (layer_0[2422] & layer_0[11174]); 
    assign out[4075] = ~(layer_0[10253] ^ layer_0[3398]); 
    assign out[4076] = ~(layer_0[218] ^ layer_0[11160]); 
    assign out[4077] = ~(layer_0[7107] & layer_0[6266]); 
    assign out[4078] = layer_0[1385] | layer_0[6242]; 
    assign out[4079] = layer_0[11210] ^ layer_0[2897]; 
    assign out[4080] = layer_0[4921] ^ layer_0[5756]; 
    assign out[4081] = layer_0[4518] ^ layer_0[8561]; 
    assign out[4082] = ~(layer_0[4546] ^ layer_0[11170]); 
    assign out[4083] = layer_0[7883] | layer_0[10689]; 
    assign out[4084] = layer_0[9928]; 
    assign out[4085] = ~layer_0[6066]; 
    assign out[4086] = ~layer_0[10682]; 
    assign out[4087] = ~(layer_0[1970] | layer_0[5712]); 
    assign out[4088] = layer_0[7018]; 
    assign out[4089] = ~layer_0[7153]; 
    assign out[4090] = layer_0[5759] ^ layer_0[6762]; 
    assign out[4091] = ~(layer_0[5154] ^ layer_0[521]); 
    assign out[4092] = ~(layer_0[3073] ^ layer_0[9502]); 
    assign out[4093] = ~(layer_0[575] | layer_0[9428]); 
    assign out[4094] = layer_0[11729] & layer_0[2573]; 
    assign out[4095] = ~(layer_0[7840] ^ layer_0[6344]); 
    assign out[4096] = ~(layer_0[9153] | layer_0[4009]); 
    assign out[4097] = layer_0[1072]; 
    assign out[4098] = layer_0[3391] ^ layer_0[5273]; 
    assign out[4099] = layer_0[3282] ^ layer_0[2649]; 
    assign out[4100] = ~layer_0[11469] | (layer_0[3180] & layer_0[11469]); 
    assign out[4101] = layer_0[4917]; 
    assign out[4102] = layer_0[9405] | layer_0[4832]; 
    assign out[4103] = layer_0[1729] ^ layer_0[932]; 
    assign out[4104] = ~(layer_0[7625] ^ layer_0[43]); 
    assign out[4105] = ~layer_0[7801] | (layer_0[7801] & layer_0[9021]); 
    assign out[4106] = ~(layer_0[3744] ^ layer_0[8698]); 
    assign out[4107] = ~layer_0[9304]; 
    assign out[4108] = ~layer_0[4634] | (layer_0[4634] & layer_0[11651]); 
    assign out[4109] = ~(layer_0[3000] & layer_0[3351]); 
    assign out[4110] = layer_0[897]; 
    assign out[4111] = ~layer_0[6243]; 
    assign out[4112] = ~(layer_0[16] ^ layer_0[5925]); 
    assign out[4113] = layer_0[1510]; 
    assign out[4114] = ~(layer_0[9924] ^ layer_0[9244]); 
    assign out[4115] = layer_0[7321] | layer_0[189]; 
    assign out[4116] = layer_0[3824] ^ layer_0[3522]; 
    assign out[4117] = layer_0[1523]; 
    assign out[4118] = ~layer_0[1859]; 
    assign out[4119] = ~(layer_0[2817] ^ layer_0[11887]); 
    assign out[4120] = ~(layer_0[7502] & layer_0[6372]); 
    assign out[4121] = ~layer_0[2671]; 
    assign out[4122] = layer_0[4757]; 
    assign out[4123] = layer_0[6394] & ~layer_0[1891]; 
    assign out[4124] = layer_0[8568]; 
    assign out[4125] = ~layer_0[5574]; 
    assign out[4126] = layer_0[1741]; 
    assign out[4127] = layer_0[5092] ^ layer_0[1570]; 
    assign out[4128] = layer_0[10590] | layer_0[6349]; 
    assign out[4129] = layer_0[7038] ^ layer_0[3986]; 
    assign out[4130] = layer_0[7851]; 
    assign out[4131] = ~layer_0[4853]; 
    assign out[4132] = ~(layer_0[9514] & layer_0[3576]); 
    assign out[4133] = layer_0[8673] & ~layer_0[9007]; 
    assign out[4134] = layer_0[11641] & layer_0[3158]; 
    assign out[4135] = layer_0[1803] & ~layer_0[8382]; 
    assign out[4136] = ~(layer_0[11779] ^ layer_0[4418]); 
    assign out[4137] = ~(layer_0[8720] ^ layer_0[4924]); 
    assign out[4138] = ~layer_0[5973]; 
    assign out[4139] = layer_0[5714] ^ layer_0[8570]; 
    assign out[4140] = ~layer_0[7437] | (layer_0[7437] & layer_0[10486]); 
    assign out[4141] = ~layer_0[5003]; 
    assign out[4142] = layer_0[1962]; 
    assign out[4143] = ~(layer_0[7050] & layer_0[6550]); 
    assign out[4144] = layer_0[10811] & layer_0[7654]; 
    assign out[4145] = ~layer_0[3615] | (layer_0[3615] & layer_0[9468]); 
    assign out[4146] = ~(layer_0[4607] ^ layer_0[846]); 
    assign out[4147] = layer_0[5011]; 
    assign out[4148] = ~(layer_0[8319] | layer_0[383]); 
    assign out[4149] = layer_0[2652]; 
    assign out[4150] = ~layer_0[6262]; 
    assign out[4151] = ~layer_0[3752]; 
    assign out[4152] = ~layer_0[6721]; 
    assign out[4153] = ~layer_0[4512] | (layer_0[4512] & layer_0[11117]); 
    assign out[4154] = ~(layer_0[2136] & layer_0[3976]); 
    assign out[4155] = layer_0[11416] | layer_0[11264]; 
    assign out[4156] = layer_0[866]; 
    assign out[4157] = ~layer_0[508]; 
    assign out[4158] = layer_0[2078] ^ layer_0[10675]; 
    assign out[4159] = ~layer_0[9427] | (layer_0[9427] & layer_0[3417]); 
    assign out[4160] = ~(layer_0[2568] ^ layer_0[10130]); 
    assign out[4161] = ~(layer_0[10182] ^ layer_0[6790]); 
    assign out[4162] = layer_0[11742]; 
    assign out[4163] = ~layer_0[4829] | (layer_0[4242] & layer_0[4829]); 
    assign out[4164] = layer_0[3089] | layer_0[2630]; 
    assign out[4165] = ~(layer_0[3221] & layer_0[10656]); 
    assign out[4166] = ~(layer_0[286] & layer_0[11289]); 
    assign out[4167] = layer_0[4447] & ~layer_0[7440]; 
    assign out[4168] = ~layer_0[4839] | (layer_0[9842] & layer_0[4839]); 
    assign out[4169] = ~layer_0[3492] | (layer_0[479] & layer_0[3492]); 
    assign out[4170] = layer_0[1708]; 
    assign out[4171] = layer_0[6065]; 
    assign out[4172] = layer_0[6733]; 
    assign out[4173] = ~layer_0[10862]; 
    assign out[4174] = layer_0[703] ^ layer_0[8970]; 
    assign out[4175] = ~(layer_0[7615] | layer_0[8974]); 
    assign out[4176] = 1'b1; 
    assign out[4177] = ~layer_0[11105] | (layer_0[11105] & layer_0[8519]); 
    assign out[4178] = layer_0[7771] & layer_0[11458]; 
    assign out[4179] = layer_0[2910]; 
    assign out[4180] = ~(layer_0[2369] ^ layer_0[11390]); 
    assign out[4181] = layer_0[10820] | layer_0[5651]; 
    assign out[4182] = ~layer_0[2475]; 
    assign out[4183] = layer_0[3503] | layer_0[3853]; 
    assign out[4184] = ~layer_0[9698] | (layer_0[9698] & layer_0[2381]); 
    assign out[4185] = layer_0[644] ^ layer_0[8923]; 
    assign out[4186] = layer_0[7675] ^ layer_0[11454]; 
    assign out[4187] = layer_0[8747] ^ layer_0[7327]; 
    assign out[4188] = ~(layer_0[6184] ^ layer_0[9718]); 
    assign out[4189] = ~(layer_0[8679] ^ layer_0[8113]); 
    assign out[4190] = layer_0[9438] ^ layer_0[11171]; 
    assign out[4191] = layer_0[9729] ^ layer_0[11041]; 
    assign out[4192] = ~(layer_0[7727] | layer_0[941]); 
    assign out[4193] = layer_0[8625]; 
    assign out[4194] = layer_0[4714] & ~layer_0[10392]; 
    assign out[4195] = ~(layer_0[2204] ^ layer_0[5576]); 
    assign out[4196] = ~layer_0[3422]; 
    assign out[4197] = ~(layer_0[2150] ^ layer_0[1407]); 
    assign out[4198] = layer_0[921]; 
    assign out[4199] = layer_0[5493]; 
    assign out[4200] = layer_0[569] | layer_0[9982]; 
    assign out[4201] = layer_0[7697] ^ layer_0[2098]; 
    assign out[4202] = ~layer_0[4038]; 
    assign out[4203] = ~(layer_0[9748] ^ layer_0[5203]); 
    assign out[4204] = layer_0[135] ^ layer_0[6016]; 
    assign out[4205] = layer_0[7653] ^ layer_0[1512]; 
    assign out[4206] = ~layer_0[4308] | (layer_0[4308] & layer_0[10093]); 
    assign out[4207] = layer_0[745] | layer_0[9913]; 
    assign out[4208] = layer_0[765] | layer_0[9634]; 
    assign out[4209] = layer_0[4616] & ~layer_0[1609]; 
    assign out[4210] = ~layer_0[7683] | (layer_0[7683] & layer_0[393]); 
    assign out[4211] = layer_0[11464] ^ layer_0[7195]; 
    assign out[4212] = ~(layer_0[766] & layer_0[7278]); 
    assign out[4213] = layer_0[1279] ^ layer_0[2740]; 
    assign out[4214] = layer_0[3259] ^ layer_0[612]; 
    assign out[4215] = layer_0[9066]; 
    assign out[4216] = layer_0[8772]; 
    assign out[4217] = ~layer_0[5046]; 
    assign out[4218] = ~layer_0[1662]; 
    assign out[4219] = layer_0[10503]; 
    assign out[4220] = layer_0[6695] & ~layer_0[268]; 
    assign out[4221] = ~(layer_0[2304] ^ layer_0[11736]); 
    assign out[4222] = ~(layer_0[8737] | layer_0[11866]); 
    assign out[4223] = layer_0[3206] | layer_0[1210]; 
    assign out[4224] = layer_0[6791] & ~layer_0[9739]; 
    assign out[4225] = layer_0[5391] ^ layer_0[5187]; 
    assign out[4226] = ~layer_0[8249]; 
    assign out[4227] = ~(layer_0[5773] | layer_0[4139]); 
    assign out[4228] = layer_0[3889] ^ layer_0[4848]; 
    assign out[4229] = layer_0[4146]; 
    assign out[4230] = layer_0[8850] & layer_0[7488]; 
    assign out[4231] = layer_0[8925] | layer_0[2917]; 
    assign out[4232] = ~layer_0[11431] | (layer_0[11431] & layer_0[2130]); 
    assign out[4233] = ~(layer_0[1389] ^ layer_0[4368]); 
    assign out[4234] = layer_0[9816]; 
    assign out[4235] = ~layer_0[5828] | (layer_0[2522] & layer_0[5828]); 
    assign out[4236] = layer_0[1086] ^ layer_0[402]; 
    assign out[4237] = layer_0[9038]; 
    assign out[4238] = layer_0[7355] & ~layer_0[1527]; 
    assign out[4239] = ~(layer_0[1192] ^ layer_0[6407]); 
    assign out[4240] = ~(layer_0[8039] | layer_0[5941]); 
    assign out[4241] = ~(layer_0[11522] & layer_0[8897]); 
    assign out[4242] = ~(layer_0[52] & layer_0[6010]); 
    assign out[4243] = ~(layer_0[9264] ^ layer_0[11930]); 
    assign out[4244] = ~layer_0[2319] | (layer_0[7260] & layer_0[2319]); 
    assign out[4245] = layer_0[1099]; 
    assign out[4246] = ~(layer_0[5114] & layer_0[6135]); 
    assign out[4247] = ~layer_0[7931]; 
    assign out[4248] = layer_0[4994]; 
    assign out[4249] = layer_0[11123] & layer_0[4846]; 
    assign out[4250] = ~(layer_0[8873] ^ layer_0[9653]); 
    assign out[4251] = layer_0[11339]; 
    assign out[4252] = layer_0[7135] ^ layer_0[9174]; 
    assign out[4253] = ~(layer_0[7539] | layer_0[833]); 
    assign out[4254] = layer_0[154]; 
    assign out[4255] = layer_0[8320]; 
    assign out[4256] = layer_0[10248] ^ layer_0[10297]; 
    assign out[4257] = layer_0[11011]; 
    assign out[4258] = layer_0[3699] & layer_0[1143]; 
    assign out[4259] = layer_0[8276] ^ layer_0[5091]; 
    assign out[4260] = ~layer_0[4750]; 
    assign out[4261] = ~(layer_0[700] ^ layer_0[5868]); 
    assign out[4262] = layer_0[4844] ^ layer_0[9185]; 
    assign out[4263] = ~(layer_0[11028] & layer_0[2139]); 
    assign out[4264] = ~layer_0[2868]; 
    assign out[4265] = ~layer_0[4750] | (layer_0[8437] & layer_0[4750]); 
    assign out[4266] = ~layer_0[3092] | (layer_0[8346] & layer_0[3092]); 
    assign out[4267] = ~layer_0[5375] | (layer_0[5375] & layer_0[1888]); 
    assign out[4268] = layer_0[2393]; 
    assign out[4269] = layer_0[7966] | layer_0[5259]; 
    assign out[4270] = ~(layer_0[536] | layer_0[8613]); 
    assign out[4271] = layer_0[6938]; 
    assign out[4272] = ~(layer_0[5446] ^ layer_0[1104]); 
    assign out[4273] = layer_0[3919] ^ layer_0[8630]; 
    assign out[4274] = ~(layer_0[1648] & layer_0[7065]); 
    assign out[4275] = ~layer_0[7120] | (layer_0[7120] & layer_0[9909]); 
    assign out[4276] = layer_0[4966] & layer_0[2834]; 
    assign out[4277] = ~(layer_0[5435] | layer_0[2325]); 
    assign out[4278] = layer_0[10635] & ~layer_0[3559]; 
    assign out[4279] = layer_0[5312] | layer_0[11125]; 
    assign out[4280] = ~layer_0[10061] | (layer_0[8678] & layer_0[10061]); 
    assign out[4281] = ~layer_0[9762]; 
    assign out[4282] = ~layer_0[9218] | (layer_0[7806] & layer_0[9218]); 
    assign out[4283] = layer_0[7616] ^ layer_0[11854]; 
    assign out[4284] = layer_0[9647]; 
    assign out[4285] = ~(layer_0[4287] ^ layer_0[45]); 
    assign out[4286] = layer_0[10555] ^ layer_0[9316]; 
    assign out[4287] = layer_0[2444] ^ layer_0[249]; 
    assign out[4288] = layer_0[11360]; 
    assign out[4289] = layer_0[2641] ^ layer_0[2460]; 
    assign out[4290] = ~layer_0[6207]; 
    assign out[4291] = layer_0[9585]; 
    assign out[4292] = ~(layer_0[1835] | layer_0[9886]); 
    assign out[4293] = ~(layer_0[5539] ^ layer_0[4537]); 
    assign out[4294] = layer_0[167]; 
    assign out[4295] = ~(layer_0[9006] | layer_0[11725]); 
    assign out[4296] = ~layer_0[8001]; 
    assign out[4297] = layer_0[9030] ^ layer_0[10735]; 
    assign out[4298] = layer_0[4803]; 
    assign out[4299] = ~layer_0[10607] | (layer_0[7106] & layer_0[10607]); 
    assign out[4300] = layer_0[5] ^ layer_0[11660]; 
    assign out[4301] = layer_0[8806] ^ layer_0[10730]; 
    assign out[4302] = ~(layer_0[9378] ^ layer_0[10887]); 
    assign out[4303] = layer_0[4290] ^ layer_0[11752]; 
    assign out[4304] = ~(layer_0[3462] | layer_0[3003]); 
    assign out[4305] = layer_0[3255]; 
    assign out[4306] = layer_0[5551] & ~layer_0[2533]; 
    assign out[4307] = layer_0[3654] ^ layer_0[9592]; 
    assign out[4308] = ~layer_0[2947]; 
    assign out[4309] = ~(layer_0[10586] ^ layer_0[2523]); 
    assign out[4310] = ~(layer_0[11891] ^ layer_0[3754]); 
    assign out[4311] = layer_0[5380] & layer_0[10142]; 
    assign out[4312] = layer_0[7021] ^ layer_0[1151]; 
    assign out[4313] = layer_0[9325]; 
    assign out[4314] = layer_0[9483] ^ layer_0[6393]; 
    assign out[4315] = layer_0[9145] ^ layer_0[5443]; 
    assign out[4316] = ~(layer_0[11659] & layer_0[6024]); 
    assign out[4317] = ~(layer_0[10603] ^ layer_0[4583]); 
    assign out[4318] = layer_0[11122]; 
    assign out[4319] = layer_0[5833] ^ layer_0[1599]; 
    assign out[4320] = ~layer_0[11245] | (layer_0[11245] & layer_0[3264]); 
    assign out[4321] = layer_0[9632] | layer_0[7229]; 
    assign out[4322] = ~(layer_0[3176] ^ layer_0[2364]); 
    assign out[4323] = ~(layer_0[6213] & layer_0[11427]); 
    assign out[4324] = layer_0[3545] ^ layer_0[378]; 
    assign out[4325] = ~layer_0[881]; 
    assign out[4326] = ~layer_0[10]; 
    assign out[4327] = ~(layer_0[930] ^ layer_0[1393]); 
    assign out[4328] = layer_0[4567]; 
    assign out[4329] = layer_0[1327]; 
    assign out[4330] = ~(layer_0[2597] ^ layer_0[3637]); 
    assign out[4331] = ~(layer_0[6934] ^ layer_0[1610]); 
    assign out[4332] = layer_0[5708]; 
    assign out[4333] = layer_0[4609] | layer_0[4237]; 
    assign out[4334] = ~layer_0[10434] | (layer_0[10434] & layer_0[1740]); 
    assign out[4335] = ~(layer_0[5431] & layer_0[9734]); 
    assign out[4336] = ~(layer_0[3720] ^ layer_0[177]); 
    assign out[4337] = ~(layer_0[6523] ^ layer_0[4367]); 
    assign out[4338] = ~layer_0[3544]; 
    assign out[4339] = ~(layer_0[3165] ^ layer_0[1558]); 
    assign out[4340] = layer_0[10079] & ~layer_0[11296]; 
    assign out[4341] = ~(layer_0[7579] & layer_0[9111]); 
    assign out[4342] = ~(layer_0[9579] ^ layer_0[6791]); 
    assign out[4343] = layer_0[7763]; 
    assign out[4344] = ~layer_0[8109]; 
    assign out[4345] = ~layer_0[541]; 
    assign out[4346] = layer_0[5046] ^ layer_0[7678]; 
    assign out[4347] = ~layer_0[8468]; 
    assign out[4348] = ~layer_0[7530]; 
    assign out[4349] = layer_0[2798]; 
    assign out[4350] = ~(layer_0[7787] & layer_0[7747]); 
    assign out[4351] = ~layer_0[2641]; 
    assign out[4352] = layer_0[5922]; 
    assign out[4353] = layer_0[9507] ^ layer_0[8298]; 
    assign out[4354] = ~(layer_0[5095] | layer_0[1134]); 
    assign out[4355] = layer_0[5455] & ~layer_0[251]; 
    assign out[4356] = ~layer_0[1854]; 
    assign out[4357] = layer_0[2001] & layer_0[8868]; 
    assign out[4358] = ~(layer_0[5661] & layer_0[9793]); 
    assign out[4359] = ~(layer_0[3920] & layer_0[10631]); 
    assign out[4360] = layer_0[3431] ^ layer_0[2595]; 
    assign out[4361] = ~(layer_0[9590] ^ layer_0[9128]); 
    assign out[4362] = layer_0[1863] | layer_0[10810]; 
    assign out[4363] = ~(layer_0[2612] ^ layer_0[10487]); 
    assign out[4364] = ~(layer_0[7500] & layer_0[275]); 
    assign out[4365] = layer_0[11313] & ~layer_0[1169]; 
    assign out[4366] = layer_0[5537] ^ layer_0[6171]; 
    assign out[4367] = layer_0[6679]; 
    assign out[4368] = layer_0[1142] ^ layer_0[11964]; 
    assign out[4369] = ~(layer_0[11306] | layer_0[6717]); 
    assign out[4370] = ~(layer_0[6705] ^ layer_0[9034]); 
    assign out[4371] = layer_0[1484] ^ layer_0[4091]; 
    assign out[4372] = ~layer_0[9763] | (layer_0[9673] & layer_0[9763]); 
    assign out[4373] = layer_0[334]; 
    assign out[4374] = layer_0[4425] ^ layer_0[1904]; 
    assign out[4375] = layer_0[2211]; 
    assign out[4376] = ~(layer_0[7508] ^ layer_0[157]); 
    assign out[4377] = layer_0[9938] ^ layer_0[7722]; 
    assign out[4378] = ~layer_0[11286]; 
    assign out[4379] = ~(layer_0[6427] ^ layer_0[11037]); 
    assign out[4380] = ~layer_0[1014]; 
    assign out[4381] = layer_0[3536] | layer_0[8520]; 
    assign out[4382] = ~layer_0[9758]; 
    assign out[4383] = ~layer_0[1465] | (layer_0[11211] & layer_0[1465]); 
    assign out[4384] = ~(layer_0[11361] ^ layer_0[3004]); 
    assign out[4385] = layer_0[2944]; 
    assign out[4386] = layer_0[2853] ^ layer_0[4332]; 
    assign out[4387] = layer_0[5772] ^ layer_0[4068]; 
    assign out[4388] = ~(layer_0[9188] & layer_0[9048]); 
    assign out[4389] = layer_0[3734] | layer_0[8456]; 
    assign out[4390] = ~layer_0[11734]; 
    assign out[4391] = ~(layer_0[3436] ^ layer_0[11911]); 
    assign out[4392] = layer_0[7511] ^ layer_0[9551]; 
    assign out[4393] = layer_0[3216] & ~layer_0[359]; 
    assign out[4394] = ~layer_0[5698]; 
    assign out[4395] = ~layer_0[7461] | (layer_0[7461] & layer_0[4883]); 
    assign out[4396] = ~(layer_0[7328] ^ layer_0[6425]); 
    assign out[4397] = ~layer_0[4359]; 
    assign out[4398] = ~layer_0[5030]; 
    assign out[4399] = layer_0[2177] & ~layer_0[17]; 
    assign out[4400] = ~(layer_0[2539] ^ layer_0[4740]); 
    assign out[4401] = ~(layer_0[8627] | layer_0[1080]); 
    assign out[4402] = layer_0[3497]; 
    assign out[4403] = ~(layer_0[8241] ^ layer_0[1075]); 
    assign out[4404] = ~(layer_0[2890] & layer_0[4109]); 
    assign out[4405] = ~layer_0[10767] | (layer_0[10767] & layer_0[11418]); 
    assign out[4406] = ~(layer_0[6991] ^ layer_0[11099]); 
    assign out[4407] = ~layer_0[9181] | (layer_0[6122] & layer_0[9181]); 
    assign out[4408] = ~layer_0[5145]; 
    assign out[4409] = ~(layer_0[8881] ^ layer_0[3240]); 
    assign out[4410] = ~(layer_0[10458] ^ layer_0[11666]); 
    assign out[4411] = layer_0[7068] & ~layer_0[5701]; 
    assign out[4412] = layer_0[4132] ^ layer_0[333]; 
    assign out[4413] = ~(layer_0[10161] ^ layer_0[11757]); 
    assign out[4414] = layer_0[9143]; 
    assign out[4415] = layer_0[2990]; 
    assign out[4416] = ~(layer_0[2670] & layer_0[8196]); 
    assign out[4417] = ~(layer_0[5681] ^ layer_0[4499]); 
    assign out[4418] = ~(layer_0[4273] ^ layer_0[4126]); 
    assign out[4419] = layer_0[4352]; 
    assign out[4420] = layer_0[1917] & layer_0[11277]; 
    assign out[4421] = layer_0[3640] & layer_0[9033]; 
    assign out[4422] = ~(layer_0[9830] ^ layer_0[7772]); 
    assign out[4423] = ~(layer_0[917] | layer_0[2445]); 
    assign out[4424] = ~(layer_0[880] & layer_0[4676]); 
    assign out[4425] = ~(layer_0[2102] ^ layer_0[10751]); 
    assign out[4426] = layer_0[852] | layer_0[4429]; 
    assign out[4427] = layer_0[4391]; 
    assign out[4428] = layer_0[1047] & layer_0[6504]; 
    assign out[4429] = layer_0[5302] ^ layer_0[4892]; 
    assign out[4430] = ~layer_0[5598] | (layer_0[5598] & layer_0[2280]); 
    assign out[4431] = layer_0[2155]; 
    assign out[4432] = layer_0[8459] & layer_0[1896]; 
    assign out[4433] = layer_0[3997] ^ layer_0[1198]; 
    assign out[4434] = ~(layer_0[9848] ^ layer_0[1608]); 
    assign out[4435] = ~(layer_0[8095] ^ layer_0[6874]); 
    assign out[4436] = layer_0[6193] | layer_0[6341]; 
    assign out[4437] = ~(layer_0[4679] ^ layer_0[8642]); 
    assign out[4438] = ~(layer_0[6300] ^ layer_0[8374]); 
    assign out[4439] = ~layer_0[9338]; 
    assign out[4440] = layer_0[1811] ^ layer_0[2517]; 
    assign out[4441] = layer_0[4314] ^ layer_0[5861]; 
    assign out[4442] = ~(layer_0[9710] ^ layer_0[6159]); 
    assign out[4443] = ~layer_0[10628] | (layer_0[10628] & layer_0[8119]); 
    assign out[4444] = layer_0[2394]; 
    assign out[4445] = layer_0[6553] & ~layer_0[4739]; 
    assign out[4446] = layer_0[8710] ^ layer_0[9080]; 
    assign out[4447] = ~(layer_0[4345] ^ layer_0[7334]); 
    assign out[4448] = ~layer_0[988] | (layer_0[988] & layer_0[9782]); 
    assign out[4449] = layer_0[8624] ^ layer_0[9810]; 
    assign out[4450] = ~layer_0[11215] | (layer_0[11215] & layer_0[5565]); 
    assign out[4451] = layer_0[1123]; 
    assign out[4452] = layer_0[11477] ^ layer_0[3093]; 
    assign out[4453] = ~layer_0[709]; 
    assign out[4454] = layer_0[8101] ^ layer_0[7251]; 
    assign out[4455] = layer_0[8243]; 
    assign out[4456] = layer_0[1093]; 
    assign out[4457] = layer_0[5578] & layer_0[2733]; 
    assign out[4458] = layer_0[6605] ^ layer_0[7632]; 
    assign out[4459] = ~layer_0[1666]; 
    assign out[4460] = layer_0[5320]; 
    assign out[4461] = ~(layer_0[7867] | layer_0[9767]); 
    assign out[4462] = ~(layer_0[9490] ^ layer_0[3914]); 
    assign out[4463] = ~layer_0[572]; 
    assign out[4464] = ~(layer_0[9556] ^ layer_0[10137]); 
    assign out[4465] = ~layer_0[11170] | (layer_0[11170] & layer_0[8889]); 
    assign out[4466] = ~layer_0[9413]; 
    assign out[4467] = layer_0[7191]; 
    assign out[4468] = layer_0[1053] ^ layer_0[456]; 
    assign out[4469] = ~layer_0[10834] | (layer_0[10834] & layer_0[4646]); 
    assign out[4470] = layer_0[7794]; 
    assign out[4471] = ~(layer_0[3814] ^ layer_0[3242]); 
    assign out[4472] = layer_0[3041]; 
    assign out[4473] = layer_0[2777] | layer_0[305]; 
    assign out[4474] = layer_0[314]; 
    assign out[4475] = layer_0[10424]; 
    assign out[4476] = ~(layer_0[6717] | layer_0[2512]); 
    assign out[4477] = layer_0[3258] | layer_0[956]; 
    assign out[4478] = ~(layer_0[11604] ^ layer_0[4903]); 
    assign out[4479] = ~(layer_0[7672] ^ layer_0[4452]); 
    assign out[4480] = ~layer_0[11860] | (layer_0[11860] & layer_0[4822]); 
    assign out[4481] = layer_0[5534] ^ layer_0[5000]; 
    assign out[4482] = layer_0[3421]; 
    assign out[4483] = layer_0[1023]; 
    assign out[4484] = layer_0[6043] & ~layer_0[6454]; 
    assign out[4485] = layer_0[8968]; 
    assign out[4486] = ~layer_0[8068]; 
    assign out[4487] = ~layer_0[2259] | (layer_0[395] & layer_0[2259]); 
    assign out[4488] = layer_0[7893] & ~layer_0[6168]; 
    assign out[4489] = layer_0[234] & ~layer_0[843]; 
    assign out[4490] = ~layer_0[2912]; 
    assign out[4491] = ~(layer_0[6507] ^ layer_0[10873]); 
    assign out[4492] = layer_0[7296] | layer_0[953]; 
    assign out[4493] = layer_0[4019] | layer_0[2604]; 
    assign out[4494] = layer_0[53] ^ layer_0[5351]; 
    assign out[4495] = ~(layer_0[11958] | layer_0[7395]); 
    assign out[4496] = layer_0[7239]; 
    assign out[4497] = ~(layer_0[7065] ^ layer_0[9508]); 
    assign out[4498] = layer_0[11592]; 
    assign out[4499] = ~layer_0[6829]; 
    assign out[4500] = ~layer_0[8184]; 
    assign out[4501] = layer_0[4017]; 
    assign out[4502] = layer_0[3338]; 
    assign out[4503] = ~layer_0[11349]; 
    assign out[4504] = layer_0[3249]; 
    assign out[4505] = layer_0[10308]; 
    assign out[4506] = ~layer_0[9841] | (layer_0[7898] & layer_0[9841]); 
    assign out[4507] = layer_0[868] ^ layer_0[5041]; 
    assign out[4508] = ~(layer_0[11478] ^ layer_0[4703]); 
    assign out[4509] = ~layer_0[7643]; 
    assign out[4510] = layer_0[9685]; 
    assign out[4511] = ~layer_0[7000]; 
    assign out[4512] = layer_0[8461] | layer_0[6123]; 
    assign out[4513] = ~layer_0[3205] | (layer_0[3205] & layer_0[6733]); 
    assign out[4514] = layer_0[316]; 
    assign out[4515] = layer_0[809] & layer_0[7902]; 
    assign out[4516] = layer_0[10555] ^ layer_0[503]; 
    assign out[4517] = layer_0[2451]; 
    assign out[4518] = ~(layer_0[10725] | layer_0[5967]); 
    assign out[4519] = ~layer_0[1515]; 
    assign out[4520] = ~layer_0[2499] | (layer_0[2499] & layer_0[5177]); 
    assign out[4521] = layer_0[10002] ^ layer_0[7446]; 
    assign out[4522] = ~(layer_0[4292] & layer_0[7289]); 
    assign out[4523] = layer_0[10273] & ~layer_0[11937]; 
    assign out[4524] = layer_0[1785] | layer_0[2102]; 
    assign out[4525] = layer_0[2962]; 
    assign out[4526] = ~(layer_0[11710] ^ layer_0[5206]); 
    assign out[4527] = layer_0[5159] ^ layer_0[515]; 
    assign out[4528] = layer_0[5724] ^ layer_0[4378]; 
    assign out[4529] = ~layer_0[550] | (layer_0[112] & layer_0[550]); 
    assign out[4530] = layer_0[4748] & ~layer_0[1839]; 
    assign out[4531] = layer_0[6492] & ~layer_0[9270]; 
    assign out[4532] = ~(layer_0[9694] ^ layer_0[10538]); 
    assign out[4533] = ~(layer_0[10621] & layer_0[2823]); 
    assign out[4534] = layer_0[6419] ^ layer_0[8359]; 
    assign out[4535] = ~layer_0[10470]; 
    assign out[4536] = layer_0[9625]; 
    assign out[4537] = ~(layer_0[3655] & layer_0[1653]); 
    assign out[4538] = layer_0[10196] ^ layer_0[11098]; 
    assign out[4539] = ~layer_0[4709] | (layer_0[4709] & layer_0[9631]); 
    assign out[4540] = layer_0[1204] | layer_0[8901]; 
    assign out[4541] = ~layer_0[2145] | (layer_0[8866] & layer_0[2145]); 
    assign out[4542] = ~(layer_0[8501] ^ layer_0[3054]); 
    assign out[4543] = layer_0[1338]; 
    assign out[4544] = ~(layer_0[1853] | layer_0[2921]); 
    assign out[4545] = layer_0[2914] & layer_0[11505]; 
    assign out[4546] = ~layer_0[1743]; 
    assign out[4547] = layer_0[9433] & ~layer_0[10797]; 
    assign out[4548] = layer_0[8404] ^ layer_0[10004]; 
    assign out[4549] = layer_0[2064]; 
    assign out[4550] = layer_0[5218] ^ layer_0[4349]; 
    assign out[4551] = ~layer_0[9173]; 
    assign out[4552] = ~layer_0[4448]; 
    assign out[4553] = ~layer_0[5886] | (layer_0[5886] & layer_0[2123]); 
    assign out[4554] = ~layer_0[6396]; 
    assign out[4555] = ~(layer_0[6437] ^ layer_0[11816]); 
    assign out[4556] = layer_0[4434]; 
    assign out[4557] = layer_0[1404] ^ layer_0[6860]; 
    assign out[4558] = ~layer_0[8830] | (layer_0[6723] & layer_0[8830]); 
    assign out[4559] = ~(layer_0[3458] ^ layer_0[11528]); 
    assign out[4560] = ~layer_0[3029]; 
    assign out[4561] = layer_0[2182] ^ layer_0[9034]; 
    assign out[4562] = ~(layer_0[737] & layer_0[2461]); 
    assign out[4563] = ~(layer_0[10466] ^ layer_0[10770]); 
    assign out[4564] = ~(layer_0[3667] & layer_0[4971]); 
    assign out[4565] = ~layer_0[2744] | (layer_0[2744] & layer_0[9566]); 
    assign out[4566] = ~(layer_0[1721] ^ layer_0[1282]); 
    assign out[4567] = ~(layer_0[4536] ^ layer_0[9363]); 
    assign out[4568] = ~(layer_0[5073] ^ layer_0[8644]); 
    assign out[4569] = ~(layer_0[5131] | layer_0[1439]); 
    assign out[4570] = ~(layer_0[5201] ^ layer_0[3439]); 
    assign out[4571] = layer_0[3070]; 
    assign out[4572] = ~layer_0[30]; 
    assign out[4573] = ~(layer_0[2342] ^ layer_0[11160]); 
    assign out[4574] = layer_0[618] | layer_0[9159]; 
    assign out[4575] = layer_0[4147]; 
    assign out[4576] = layer_0[1914] ^ layer_0[9615]; 
    assign out[4577] = layer_0[9369] | layer_0[813]; 
    assign out[4578] = layer_0[3549]; 
    assign out[4579] = layer_0[4228] ^ layer_0[9118]; 
    assign out[4580] = layer_0[7425] & layer_0[112]; 
    assign out[4581] = layer_0[2174] & ~layer_0[2699]; 
    assign out[4582] = layer_0[11546] ^ layer_0[4756]; 
    assign out[4583] = ~(layer_0[426] ^ layer_0[9701]); 
    assign out[4584] = ~(layer_0[10508] ^ layer_0[1828]); 
    assign out[4585] = layer_0[450]; 
    assign out[4586] = ~(layer_0[2647] ^ layer_0[9775]); 
    assign out[4587] = ~(layer_0[815] & layer_0[872]); 
    assign out[4588] = ~layer_0[9961]; 
    assign out[4589] = layer_0[10011] & layer_0[3403]; 
    assign out[4590] = ~layer_0[5386]; 
    assign out[4591] = ~(layer_0[11026] ^ layer_0[2774]); 
    assign out[4592] = layer_0[6529]; 
    assign out[4593] = layer_0[11811] | layer_0[9795]; 
    assign out[4594] = layer_0[6575] & ~layer_0[11506]; 
    assign out[4595] = layer_0[696]; 
    assign out[4596] = ~(layer_0[5369] ^ layer_0[10915]); 
    assign out[4597] = ~(layer_0[3226] ^ layer_0[1756]); 
    assign out[4598] = layer_0[1538] | layer_0[1923]; 
    assign out[4599] = layer_0[6294] | layer_0[6977]; 
    assign out[4600] = ~layer_0[8315] | (layer_0[9435] & layer_0[8315]); 
    assign out[4601] = ~(layer_0[9970] | layer_0[5477]); 
    assign out[4602] = layer_0[1416] | layer_0[3363]; 
    assign out[4603] = ~layer_0[11374] | (layer_0[2505] & layer_0[11374]); 
    assign out[4604] = ~layer_0[9060]; 
    assign out[4605] = ~(layer_0[9637] ^ layer_0[1137]); 
    assign out[4606] = ~(layer_0[7889] ^ layer_0[6197]); 
    assign out[4607] = ~(layer_0[1095] & layer_0[485]); 
    assign out[4608] = ~layer_0[3433] | (layer_0[10968] & layer_0[3433]); 
    assign out[4609] = ~layer_0[2906]; 
    assign out[4610] = ~layer_0[7104]; 
    assign out[4611] = ~(layer_0[11204] ^ layer_0[8971]); 
    assign out[4612] = ~(layer_0[3941] ^ layer_0[8758]); 
    assign out[4613] = ~layer_0[6627]; 
    assign out[4614] = layer_0[5347] ^ layer_0[4771]; 
    assign out[4615] = layer_0[7222] ^ layer_0[6340]; 
    assign out[4616] = ~(layer_0[6040] ^ layer_0[4591]); 
    assign out[4617] = ~layer_0[7292] | (layer_0[11082] & layer_0[7292]); 
    assign out[4618] = ~layer_0[4461]; 
    assign out[4619] = ~layer_0[5326]; 
    assign out[4620] = ~(layer_0[952] & layer_0[9002]); 
    assign out[4621] = ~(layer_0[1079] | layer_0[1625]); 
    assign out[4622] = layer_0[6177] | layer_0[790]; 
    assign out[4623] = ~layer_0[4913]; 
    assign out[4624] = layer_0[9488]; 
    assign out[4625] = layer_0[2030] ^ layer_0[5769]; 
    assign out[4626] = ~layer_0[2285]; 
    assign out[4627] = 1'b1; 
    assign out[4628] = ~(layer_0[3085] | layer_0[2502]); 
    assign out[4629] = layer_0[6368] ^ layer_0[10037]; 
    assign out[4630] = ~(layer_0[10520] ^ layer_0[1266]); 
    assign out[4631] = layer_0[11398]; 
    assign out[4632] = layer_0[3543] & layer_0[5023]; 
    assign out[4633] = ~(layer_0[4999] | layer_0[4054]); 
    assign out[4634] = layer_0[11525] & layer_0[11074]; 
    assign out[4635] = ~(layer_0[11971] ^ layer_0[3220]); 
    assign out[4636] = ~layer_0[10733]; 
    assign out[4637] = ~layer_0[6004] | (layer_0[6004] & layer_0[3970]); 
    assign out[4638] = ~(layer_0[1426] ^ layer_0[4806]); 
    assign out[4639] = ~layer_0[8002]; 
    assign out[4640] = ~layer_0[3106]; 
    assign out[4641] = ~layer_0[1837]; 
    assign out[4642] = layer_0[10382]; 
    assign out[4643] = layer_0[5846] & ~layer_0[6858]; 
    assign out[4644] = ~layer_0[4074]; 
    assign out[4645] = ~layer_0[7138] | (layer_0[10322] & layer_0[7138]); 
    assign out[4646] = layer_0[2506] & ~layer_0[8128]; 
    assign out[4647] = layer_0[2809] | layer_0[7449]; 
    assign out[4648] = ~layer_0[5453] | (layer_0[10507] & layer_0[5453]); 
    assign out[4649] = ~layer_0[5992] | (layer_0[3386] & layer_0[5992]); 
    assign out[4650] = layer_0[3694]; 
    assign out[4651] = ~layer_0[3408]; 
    assign out[4652] = ~layer_0[929]; 
    assign out[4653] = layer_0[8432] & ~layer_0[8771]; 
    assign out[4654] = layer_0[8282] & ~layer_0[4026]; 
    assign out[4655] = ~layer_0[5788] | (layer_0[6756] & layer_0[5788]); 
    assign out[4656] = layer_0[4937]; 
    assign out[4657] = ~layer_0[7895]; 
    assign out[4658] = ~layer_0[10866]; 
    assign out[4659] = layer_0[9975] & ~layer_0[8117]; 
    assign out[4660] = ~layer_0[6685] | (layer_0[1685] & layer_0[6685]); 
    assign out[4661] = layer_0[8622] ^ layer_0[10252]; 
    assign out[4662] = ~layer_0[11709]; 
    assign out[4663] = layer_0[5352] | layer_0[2669]; 
    assign out[4664] = ~layer_0[3382]; 
    assign out[4665] = ~layer_0[323]; 
    assign out[4666] = layer_0[7286]; 
    assign out[4667] = ~layer_0[7728] | (layer_0[7728] & layer_0[6588]); 
    assign out[4668] = ~(layer_0[3407] ^ layer_0[6697]); 
    assign out[4669] = layer_0[11409]; 
    assign out[4670] = layer_0[11434]; 
    assign out[4671] = ~layer_0[8628]; 
    assign out[4672] = layer_0[7527]; 
    assign out[4673] = ~layer_0[2199]; 
    assign out[4674] = ~(layer_0[9370] & layer_0[5390]); 
    assign out[4675] = ~layer_0[2008]; 
    assign out[4676] = layer_0[2087]; 
    assign out[4677] = layer_0[1929] ^ layer_0[8413]; 
    assign out[4678] = ~layer_0[8954] | (layer_0[8954] & layer_0[10126]); 
    assign out[4679] = layer_0[3683] ^ layer_0[11851]; 
    assign out[4680] = layer_0[8208] & layer_0[8490]; 
    assign out[4681] = layer_0[5823] | layer_0[5984]; 
    assign out[4682] = layer_0[11043] ^ layer_0[8336]; 
    assign out[4683] = ~layer_0[5954] | (layer_0[5954] & layer_0[8299]); 
    assign out[4684] = ~layer_0[337] | (layer_0[1615] & layer_0[337]); 
    assign out[4685] = layer_0[8952] ^ layer_0[803]; 
    assign out[4686] = layer_0[581] & layer_0[6766]; 
    assign out[4687] = layer_0[7277] & layer_0[6646]; 
    assign out[4688] = layer_0[9013] ^ layer_0[1364]; 
    assign out[4689] = layer_0[7821]; 
    assign out[4690] = layer_0[5776] & ~layer_0[11180]; 
    assign out[4691] = ~(layer_0[8215] & layer_0[3346]); 
    assign out[4692] = layer_0[6742] ^ layer_0[5389]; 
    assign out[4693] = layer_0[11690]; 
    assign out[4694] = layer_0[220] & ~layer_0[5114]; 
    assign out[4695] = layer_0[7062] | layer_0[3768]; 
    assign out[4696] = ~layer_0[204]; 
    assign out[4697] = layer_0[7748] ^ layer_0[6420]; 
    assign out[4698] = ~(layer_0[11466] ^ layer_0[11567]); 
    assign out[4699] = layer_0[5595] ^ layer_0[6974]; 
    assign out[4700] = layer_0[671] | layer_0[3424]; 
    assign out[4701] = layer_0[7959] ^ layer_0[10461]; 
    assign out[4702] = layer_0[938] & ~layer_0[2202]; 
    assign out[4703] = layer_0[7175]; 
    assign out[4704] = ~(layer_0[3413] ^ layer_0[3369]); 
    assign out[4705] = ~(layer_0[5762] ^ layer_0[5723]); 
    assign out[4706] = ~(layer_0[5800] ^ layer_0[6585]); 
    assign out[4707] = layer_0[6995] & layer_0[4263]; 
    assign out[4708] = layer_0[3449] & layer_0[10653]; 
    assign out[4709] = ~layer_0[1028] | (layer_0[1028] & layer_0[561]); 
    assign out[4710] = ~(layer_0[5262] | layer_0[10082]); 
    assign out[4711] = ~(layer_0[7648] ^ layer_0[313]); 
    assign out[4712] = layer_0[6736] ^ layer_0[6700]; 
    assign out[4713] = ~layer_0[11266]; 
    assign out[4714] = layer_0[5294] & ~layer_0[1848]; 
    assign out[4715] = layer_0[8585] & ~layer_0[6131]; 
    assign out[4716] = layer_0[5420] ^ layer_0[10053]; 
    assign out[4717] = ~(layer_0[7292] | layer_0[1951]); 
    assign out[4718] = layer_0[11448] | layer_0[6224]; 
    assign out[4719] = layer_0[3071] | layer_0[7197]; 
    assign out[4720] = layer_0[6332] & ~layer_0[8090]; 
    assign out[4721] = ~(layer_0[1629] & layer_0[767]); 
    assign out[4722] = ~(layer_0[2714] | layer_0[8141]); 
    assign out[4723] = layer_0[9520] & layer_0[8664]; 
    assign out[4724] = ~layer_0[394] | (layer_0[394] & layer_0[4986]); 
    assign out[4725] = ~layer_0[2524]; 
    assign out[4726] = layer_0[11077] | layer_0[11462]; 
    assign out[4727] = ~(layer_0[818] | layer_0[2648]); 
    assign out[4728] = layer_0[7116] & ~layer_0[11324]; 
    assign out[4729] = ~layer_0[1666]; 
    assign out[4730] = ~(layer_0[7020] & layer_0[5911]); 
    assign out[4731] = layer_0[1902] | layer_0[2173]; 
    assign out[4732] = ~layer_0[1658] | (layer_0[1658] & layer_0[1002]); 
    assign out[4733] = ~layer_0[278] | (layer_0[7450] & layer_0[278]); 
    assign out[4734] = ~(layer_0[6229] ^ layer_0[4692]); 
    assign out[4735] = ~layer_0[7560]; 
    assign out[4736] = layer_0[11582]; 
    assign out[4737] = ~layer_0[8079] | (layer_0[8079] & layer_0[7968]); 
    assign out[4738] = layer_0[5935]; 
    assign out[4739] = layer_0[4211]; 
    assign out[4740] = layer_0[3928]; 
    assign out[4741] = layer_0[11235] ^ layer_0[2964]; 
    assign out[4742] = layer_0[5283] & ~layer_0[7474]; 
    assign out[4743] = layer_0[10420]; 
    assign out[4744] = ~layer_0[6053]; 
    assign out[4745] = layer_0[8047] & ~layer_0[11797]; 
    assign out[4746] = ~(layer_0[166] ^ layer_0[5150]); 
    assign out[4747] = ~(layer_0[478] ^ layer_0[8702]); 
    assign out[4748] = layer_0[3557] | layer_0[4177]; 
    assign out[4749] = ~layer_0[4123] | (layer_0[4123] & layer_0[1601]); 
    assign out[4750] = layer_0[2837] ^ layer_0[5252]; 
    assign out[4751] = ~layer_0[5510] | (layer_0[6909] & layer_0[5510]); 
    assign out[4752] = layer_0[1596] & ~layer_0[4187]; 
    assign out[4753] = layer_0[6696] | layer_0[7287]; 
    assign out[4754] = layer_0[9996] ^ layer_0[3623]; 
    assign out[4755] = ~layer_0[416] | (layer_0[8447] & layer_0[416]); 
    assign out[4756] = ~(layer_0[2609] | layer_0[5519]); 
    assign out[4757] = layer_0[6126] | layer_0[5101]; 
    assign out[4758] = layer_0[7855]; 
    assign out[4759] = layer_0[10409] ^ layer_0[4725]; 
    assign out[4760] = ~layer_0[1007]; 
    assign out[4761] = ~layer_0[11424] | (layer_0[6622] & layer_0[11424]); 
    assign out[4762] = ~(layer_0[6907] ^ layer_0[9536]); 
    assign out[4763] = ~layer_0[10346] | (layer_0[10346] & layer_0[10869]); 
    assign out[4764] = layer_0[1009] | layer_0[8302]; 
    assign out[4765] = ~layer_0[2492] | (layer_0[11894] & layer_0[2492]); 
    assign out[4766] = layer_0[11246] ^ layer_0[639]; 
    assign out[4767] = ~layer_0[2249]; 
    assign out[4768] = layer_0[11410] ^ layer_0[8010]; 
    assign out[4769] = layer_0[4375] & ~layer_0[11684]; 
    assign out[4770] = layer_0[1423]; 
    assign out[4771] = ~(layer_0[7010] & layer_0[201]); 
    assign out[4772] = layer_0[7069] ^ layer_0[1341]; 
    assign out[4773] = layer_0[8723] | layer_0[1983]; 
    assign out[4774] = layer_0[7829] ^ layer_0[2075]; 
    assign out[4775] = layer_0[7674]; 
    assign out[4776] = ~(layer_0[7138] ^ layer_0[11589]); 
    assign out[4777] = layer_0[11645] ^ layer_0[6451]; 
    assign out[4778] = ~layer_0[4988]; 
    assign out[4779] = ~(layer_0[8576] & layer_0[1668]); 
    assign out[4780] = layer_0[11188]; 
    assign out[4781] = ~layer_0[958]; 
    assign out[4782] = layer_0[7947] ^ layer_0[2599]; 
    assign out[4783] = ~(layer_0[7566] ^ layer_0[1199]); 
    assign out[4784] = layer_0[3949] ^ layer_0[1628]; 
    assign out[4785] = layer_0[5282]; 
    assign out[4786] = layer_0[9589]; 
    assign out[4787] = layer_0[531]; 
    assign out[4788] = ~(layer_0[10314] & layer_0[5556]); 
    assign out[4789] = ~(layer_0[6574] & layer_0[1990]); 
    assign out[4790] = ~layer_0[5556] | (layer_0[11452] & layer_0[5556]); 
    assign out[4791] = layer_0[7112]; 
    assign out[4792] = layer_0[7641] ^ layer_0[8982]; 
    assign out[4793] = layer_0[7924]; 
    assign out[4794] = ~layer_0[4348]; 
    assign out[4795] = layer_0[9394]; 
    assign out[4796] = ~layer_0[11616] | (layer_0[11616] & layer_0[2977]); 
    assign out[4797] = layer_0[11716] ^ layer_0[1026]; 
    assign out[4798] = ~layer_0[10611] | (layer_0[10611] & layer_0[2704]); 
    assign out[4799] = ~layer_0[2446]; 
    assign out[4800] = layer_0[7181] & ~layer_0[5036]; 
    assign out[4801] = layer_0[7863] | layer_0[1933]; 
    assign out[4802] = layer_0[10127]; 
    assign out[4803] = layer_0[11811] ^ layer_0[9090]; 
    assign out[4804] = ~(layer_0[3654] ^ layer_0[6546]); 
    assign out[4805] = layer_0[6]; 
    assign out[4806] = layer_0[10452]; 
    assign out[4807] = ~(layer_0[537] ^ layer_0[11958]); 
    assign out[4808] = ~(layer_0[1831] & layer_0[4585]); 
    assign out[4809] = layer_0[10114] ^ layer_0[4118]; 
    assign out[4810] = ~(layer_0[8864] ^ layer_0[7817]); 
    assign out[4811] = ~(layer_0[4731] ^ layer_0[9382]); 
    assign out[4812] = ~(layer_0[176] ^ layer_0[4318]); 
    assign out[4813] = ~(layer_0[9788] ^ layer_0[8235]); 
    assign out[4814] = layer_0[9732] ^ layer_0[10070]; 
    assign out[4815] = ~(layer_0[10568] | layer_0[2036]); 
    assign out[4816] = layer_0[3905] & ~layer_0[1718]; 
    assign out[4817] = layer_0[317] & ~layer_0[1354]; 
    assign out[4818] = layer_0[321] ^ layer_0[2506]; 
    assign out[4819] = layer_0[9860] ^ layer_0[824]; 
    assign out[4820] = layer_0[6003] ^ layer_0[9068]; 
    assign out[4821] = ~(layer_0[5336] & layer_0[5108]); 
    assign out[4822] = ~layer_0[7160]; 
    assign out[4823] = ~(layer_0[2140] ^ layer_0[7836]); 
    assign out[4824] = layer_0[5782] & ~layer_0[11323]; 
    assign out[4825] = layer_0[8395] | layer_0[730]; 
    assign out[4826] = ~(layer_0[10922] & layer_0[3173]); 
    assign out[4827] = layer_0[9146] ^ layer_0[6700]; 
    assign out[4828] = layer_0[9798] ^ layer_0[368]; 
    assign out[4829] = layer_0[8427] ^ layer_0[972]; 
    assign out[4830] = layer_0[11126]; 
    assign out[4831] = layer_0[7250] ^ layer_0[4768]; 
    assign out[4832] = layer_0[11252] ^ layer_0[738]; 
    assign out[4833] = ~(layer_0[3322] ^ layer_0[8158]); 
    assign out[4834] = ~(layer_0[4941] ^ layer_0[10604]); 
    assign out[4835] = layer_0[7946]; 
    assign out[4836] = layer_0[3074] & ~layer_0[2397]; 
    assign out[4837] = layer_0[10691] ^ layer_0[9569]; 
    assign out[4838] = layer_0[1980] ^ layer_0[589]; 
    assign out[4839] = ~layer_0[692]; 
    assign out[4840] = ~layer_0[5900]; 
    assign out[4841] = ~(layer_0[5695] ^ layer_0[6792]); 
    assign out[4842] = ~(layer_0[3530] ^ layer_0[10519]); 
    assign out[4843] = ~layer_0[7614] | (layer_0[1531] & layer_0[7614]); 
    assign out[4844] = ~(layer_0[6804] ^ layer_0[905]); 
    assign out[4845] = layer_0[10486] ^ layer_0[5395]; 
    assign out[4846] = layer_0[10218] & layer_0[3939]; 
    assign out[4847] = layer_0[7603] & ~layer_0[4551]; 
    assign out[4848] = layer_0[645] & ~layer_0[8200]; 
    assign out[4849] = ~(layer_0[9505] ^ layer_0[11980]); 
    assign out[4850] = ~(layer_0[7751] & layer_0[4981]); 
    assign out[4851] = ~(layer_0[10680] ^ layer_0[9456]); 
    assign out[4852] = layer_0[9169] ^ layer_0[4326]; 
    assign out[4853] = ~(layer_0[2215] | layer_0[11644]); 
    assign out[4854] = ~(layer_0[6558] ^ layer_0[1122]); 
    assign out[4855] = layer_0[2583] ^ layer_0[4736]; 
    assign out[4856] = layer_0[5874] & ~layer_0[5880]; 
    assign out[4857] = ~layer_0[9255] | (layer_0[3666] & layer_0[9255]); 
    assign out[4858] = ~(layer_0[4888] ^ layer_0[7948]); 
    assign out[4859] = layer_0[9009] & layer_0[3134]; 
    assign out[4860] = ~(layer_0[4753] ^ layer_0[687]); 
    assign out[4861] = layer_0[10678] & ~layer_0[1391]; 
    assign out[4862] = layer_0[2183] ^ layer_0[8322]; 
    assign out[4863] = layer_0[3077] ^ layer_0[5792]; 
    assign out[4864] = ~(layer_0[1247] ^ layer_0[211]); 
    assign out[4865] = ~(layer_0[6460] ^ layer_0[3028]); 
    assign out[4866] = layer_0[3138] ^ layer_0[912]; 
    assign out[4867] = ~(layer_0[10638] ^ layer_0[11565]); 
    assign out[4868] = ~(layer_0[8962] ^ layer_0[4515]); 
    assign out[4869] = layer_0[11148] ^ layer_0[10706]; 
    assign out[4870] = ~(layer_0[8347] ^ layer_0[5583]); 
    assign out[4871] = ~(layer_0[11642] ^ layer_0[5222]); 
    assign out[4872] = ~layer_0[1676]; 
    assign out[4873] = layer_0[10948]; 
    assign out[4874] = layer_0[7956]; 
    assign out[4875] = layer_0[2469] ^ layer_0[7283]; 
    assign out[4876] = layer_0[10283]; 
    assign out[4877] = layer_0[5545] & layer_0[8021]; 
    assign out[4878] = ~layer_0[3899] | (layer_0[9216] & layer_0[3899]); 
    assign out[4879] = layer_0[9352] ^ layer_0[11467]; 
    assign out[4880] = ~(layer_0[436] ^ layer_0[9720]); 
    assign out[4881] = layer_0[9138]; 
    assign out[4882] = ~(layer_0[7861] ^ layer_0[1877]); 
    assign out[4883] = layer_0[2338] ^ layer_0[7505]; 
    assign out[4884] = layer_0[10081]; 
    assign out[4885] = ~(layer_0[1491] ^ layer_0[4485]); 
    assign out[4886] = layer_0[4112] ^ layer_0[10904]; 
    assign out[4887] = layer_0[10221]; 
    assign out[4888] = ~(layer_0[7465] ^ layer_0[2653]); 
    assign out[4889] = ~(layer_0[6817] ^ layer_0[4495]); 
    assign out[4890] = layer_0[47] ^ layer_0[8000]; 
    assign out[4891] = layer_0[4732] ^ layer_0[668]; 
    assign out[4892] = layer_0[538] ^ layer_0[8095]; 
    assign out[4893] = ~layer_0[1586]; 
    assign out[4894] = ~(layer_0[326] & layer_0[1907]); 
    assign out[4895] = ~layer_0[11893] | (layer_0[3497] & layer_0[11893]); 
    assign out[4896] = layer_0[7883] | layer_0[10918]; 
    assign out[4897] = ~(layer_0[3428] ^ layer_0[8132]); 
    assign out[4898] = ~layer_0[9080] | (layer_0[9080] & layer_0[3588]); 
    assign out[4899] = ~(layer_0[8212] ^ layer_0[7516]); 
    assign out[4900] = ~layer_0[9636]; 
    assign out[4901] = ~(layer_0[969] ^ layer_0[10449]); 
    assign out[4902] = ~(layer_0[10604] ^ layer_0[2608]); 
    assign out[4903] = layer_0[3535] ^ layer_0[6333]; 
    assign out[4904] = layer_0[424] | layer_0[10263]; 
    assign out[4905] = ~(layer_0[981] & layer_0[6619]); 
    assign out[4906] = ~(layer_0[1083] & layer_0[10110]); 
    assign out[4907] = layer_0[9769] ^ layer_0[2540]; 
    assign out[4908] = ~(layer_0[2254] | layer_0[11929]); 
    assign out[4909] = ~(layer_0[10774] ^ layer_0[7499]); 
    assign out[4910] = ~layer_0[8259] | (layer_0[10654] & layer_0[8259]); 
    assign out[4911] = layer_0[3542] & ~layer_0[50]; 
    assign out[4912] = ~layer_0[7844]; 
    assign out[4913] = ~(layer_0[1339] & layer_0[9756]); 
    assign out[4914] = ~layer_0[354] | (layer_0[10794] & layer_0[354]); 
    assign out[4915] = ~layer_0[3246]; 
    assign out[4916] = ~(layer_0[10598] & layer_0[11740]); 
    assign out[4917] = layer_0[7227] ^ layer_0[5343]; 
    assign out[4918] = ~(layer_0[10618] ^ layer_0[3268]); 
    assign out[4919] = ~(layer_0[4914] ^ layer_0[7209]); 
    assign out[4920] = ~layer_0[11016]; 
    assign out[4921] = layer_0[7009] & ~layer_0[2174]; 
    assign out[4922] = layer_0[7686] ^ layer_0[9119]; 
    assign out[4923] = ~layer_0[3993]; 
    assign out[4924] = layer_0[4730] ^ layer_0[11197]; 
    assign out[4925] = layer_0[798] ^ layer_0[11873]; 
    assign out[4926] = layer_0[9236] ^ layer_0[6094]; 
    assign out[4927] = layer_0[7169]; 
    assign out[4928] = layer_0[4868] ^ layer_0[4270]; 
    assign out[4929] = ~(layer_0[11485] ^ layer_0[6328]); 
    assign out[4930] = layer_0[8364] ^ layer_0[7788]; 
    assign out[4931] = layer_0[4430] | layer_0[2950]; 
    assign out[4932] = ~(layer_0[2935] ^ layer_0[2066]); 
    assign out[4933] = layer_0[720] & ~layer_0[11987]; 
    assign out[4934] = ~(layer_0[7923] | layer_0[2560]); 
    assign out[4935] = layer_0[10399] ^ layer_0[3579]; 
    assign out[4936] = ~(layer_0[193] ^ layer_0[4612]); 
    assign out[4937] = ~(layer_0[2716] ^ layer_0[9621]); 
    assign out[4938] = ~layer_0[8073]; 
    assign out[4939] = layer_0[4857] | layer_0[5055]; 
    assign out[4940] = layer_0[5621] ^ layer_0[8852]; 
    assign out[4941] = layer_0[7157] ^ layer_0[7905]; 
    assign out[4942] = layer_0[9056] & layer_0[1114]; 
    assign out[4943] = ~(layer_0[459] ^ layer_0[11356]); 
    assign out[4944] = ~(layer_0[7988] ^ layer_0[1585]); 
    assign out[4945] = layer_0[2265] & layer_0[5954]; 
    assign out[4946] = layer_0[6871]; 
    assign out[4947] = layer_0[3281] ^ layer_0[10975]; 
    assign out[4948] = layer_0[11791] & ~layer_0[5881]; 
    assign out[4949] = layer_0[5647] ^ layer_0[6411]; 
    assign out[4950] = ~(layer_0[2438] ^ layer_0[3770]); 
    assign out[4951] = ~(layer_0[11807] ^ layer_0[5077]); 
    assign out[4952] = ~(layer_0[3991] | layer_0[8795]); 
    assign out[4953] = ~(layer_0[6215] ^ layer_0[7099]); 
    assign out[4954] = layer_0[3968] | layer_0[1105]; 
    assign out[4955] = layer_0[2086] ^ layer_0[1184]; 
    assign out[4956] = ~(layer_0[2925] ^ layer_0[7541]); 
    assign out[4957] = ~(layer_0[9721] | layer_0[174]); 
    assign out[4958] = ~(layer_0[4980] & layer_0[4463]); 
    assign out[4959] = ~(layer_0[10391] ^ layer_0[4629]); 
    assign out[4960] = layer_0[1223]; 
    assign out[4961] = ~layer_0[7888]; 
    assign out[4962] = ~layer_0[4364]; 
    assign out[4963] = ~(layer_0[1064] | layer_0[10073]); 
    assign out[4964] = ~(layer_0[1030] | layer_0[5600]); 
    assign out[4965] = layer_0[995]; 
    assign out[4966] = ~(layer_0[2374] ^ layer_0[2067]); 
    assign out[4967] = ~(layer_0[9845] | layer_0[11839]); 
    assign out[4968] = ~(layer_0[1328] ^ layer_0[2044]); 
    assign out[4969] = layer_0[10169] ^ layer_0[2667]; 
    assign out[4970] = ~(layer_0[4620] ^ layer_0[8049]); 
    assign out[4971] = ~(layer_0[3448] & layer_0[4234]); 
    assign out[4972] = ~(layer_0[324] & layer_0[6116]); 
    assign out[4973] = ~(layer_0[5020] ^ layer_0[11634]); 
    assign out[4974] = ~(layer_0[10014] ^ layer_0[11885]); 
    assign out[4975] = layer_0[7572] ^ layer_0[9301]; 
    assign out[4976] = layer_0[3629] & layer_0[5213]; 
    assign out[4977] = layer_0[7864] ^ layer_0[5789]; 
    assign out[4978] = ~layer_0[8495] | (layer_0[8495] & layer_0[7816]); 
    assign out[4979] = ~(layer_0[1508] ^ layer_0[5836]); 
    assign out[4980] = layer_0[9055] ^ layer_0[724]; 
    assign out[4981] = layer_0[5639] ^ layer_0[6989]; 
    assign out[4982] = ~layer_0[657]; 
    assign out[4983] = ~layer_0[6818]; 
    assign out[4984] = ~layer_0[9949]; 
    assign out[4985] = layer_0[6145] | layer_0[10868]; 
    assign out[4986] = layer_0[3440] & ~layer_0[9808]; 
    assign out[4987] = ~layer_0[11028]; 
    assign out[4988] = layer_0[3677]; 
    assign out[4989] = ~(layer_0[10894] ^ layer_0[7766]); 
    assign out[4990] = layer_0[10398] | layer_0[4336]; 
    assign out[4991] = ~layer_0[2352] | (layer_0[1714] & layer_0[2352]); 
    assign out[4992] = ~layer_0[9811]; 
    assign out[4993] = ~(layer_0[5134] ^ layer_0[10351]); 
    assign out[4994] = layer_0[6878] & ~layer_0[2805]; 
    assign out[4995] = ~(layer_0[3370] | layer_0[169]); 
    assign out[4996] = ~(layer_0[10171] ^ layer_0[8123]); 
    assign out[4997] = ~layer_0[9865] | (layer_0[9865] & layer_0[9862]); 
    assign out[4998] = layer_0[8135] ^ layer_0[7032]; 
    assign out[4999] = ~layer_0[991]; 
    assign out[5000] = ~(layer_0[11422] ^ layer_0[9999]); 
    assign out[5001] = layer_0[5058] ^ layer_0[3179]; 
    assign out[5002] = layer_0[6601] & ~layer_0[1983]; 
    assign out[5003] = layer_0[124] ^ layer_0[1566]; 
    assign out[5004] = ~(layer_0[11306] ^ layer_0[3395]); 
    assign out[5005] = ~layer_0[4548]; 
    assign out[5006] = layer_0[6335] ^ layer_0[790]; 
    assign out[5007] = layer_0[2482] ^ layer_0[11267]; 
    assign out[5008] = ~(layer_0[3360] & layer_0[10455]); 
    assign out[5009] = ~layer_0[2039]; 
    assign out[5010] = ~layer_0[7935] | (layer_0[3573] & layer_0[7935]); 
    assign out[5011] = ~(layer_0[8225] ^ layer_0[1258]); 
    assign out[5012] = layer_0[6447] ^ layer_0[8924]; 
    assign out[5013] = ~(layer_0[2653] ^ layer_0[4409]); 
    assign out[5014] = layer_0[5221] | layer_0[878]; 
    assign out[5015] = ~layer_0[5152] | (layer_0[697] & layer_0[5152]); 
    assign out[5016] = ~(layer_0[9276] & layer_0[11512]); 
    assign out[5017] = layer_0[10997] ^ layer_0[5125]; 
    assign out[5018] = layer_0[4591] & layer_0[1934]; 
    assign out[5019] = layer_0[8726]; 
    assign out[5020] = ~(layer_0[10729] ^ layer_0[6029]); 
    assign out[5021] = ~(layer_0[8695] ^ layer_0[1071]); 
    assign out[5022] = ~(layer_0[5694] ^ layer_0[5293]); 
    assign out[5023] = layer_0[8960]; 
    assign out[5024] = ~(layer_0[4122] ^ layer_0[5261]); 
    assign out[5025] = layer_0[5678] ^ layer_0[3058]; 
    assign out[5026] = layer_0[5978] ^ layer_0[512]; 
    assign out[5027] = ~(layer_0[7459] ^ layer_0[5025]); 
    assign out[5028] = layer_0[1988] ^ layer_0[7396]; 
    assign out[5029] = ~(layer_0[11231] & layer_0[10742]); 
    assign out[5030] = ~(layer_0[11300] ^ layer_0[1305]); 
    assign out[5031] = layer_0[4911] ^ layer_0[10453]; 
    assign out[5032] = ~(layer_0[2106] ^ layer_0[2556]); 
    assign out[5033] = layer_0[1399] & layer_0[11346]; 
    assign out[5034] = ~layer_0[11538]; 
    assign out[5035] = ~layer_0[9025]; 
    assign out[5036] = ~(layer_0[1806] | layer_0[2585]); 
    assign out[5037] = layer_0[1921] ^ layer_0[7123]; 
    assign out[5038] = ~(layer_0[1246] ^ layer_0[10092]); 
    assign out[5039] = ~(layer_0[5671] ^ layer_0[6628]); 
    assign out[5040] = layer_0[10558] & ~layer_0[10769]; 
    assign out[5041] = ~(layer_0[2731] & layer_0[9243]); 
    assign out[5042] = ~layer_0[7497]; 
    assign out[5043] = ~(layer_0[3117] ^ layer_0[11731]); 
    assign out[5044] = layer_0[4439] & ~layer_0[9834]; 
    assign out[5045] = layer_0[7071] ^ layer_0[8130]; 
    assign out[5046] = layer_0[5598] & ~layer_0[2515]; 
    assign out[5047] = layer_0[1257] ^ layer_0[2278]; 
    assign out[5048] = layer_0[7336] | layer_0[9551]; 
    assign out[5049] = ~(layer_0[3362] ^ layer_0[8439]); 
    assign out[5050] = layer_0[11412] ^ layer_0[4299]; 
    assign out[5051] = ~(layer_0[2886] ^ layer_0[8439]); 
    assign out[5052] = ~(layer_0[4274] ^ layer_0[2745]); 
    assign out[5053] = layer_0[7077]; 
    assign out[5054] = ~layer_0[6796]; 
    assign out[5055] = ~(layer_0[10329] ^ layer_0[8436]); 
    assign out[5056] = layer_0[1330] & ~layer_0[11465]; 
    assign out[5057] = ~(layer_0[3237] ^ layer_0[8087]); 
    assign out[5058] = layer_0[11202] ^ layer_0[6187]; 
    assign out[5059] = ~layer_0[2306]; 
    assign out[5060] = ~(layer_0[7384] ^ layer_0[4835]); 
    assign out[5061] = ~layer_0[6217]; 
    assign out[5062] = ~(layer_0[10698] ^ layer_0[6023]); 
    assign out[5063] = layer_0[11417]; 
    assign out[5064] = ~layer_0[10963] | (layer_0[10963] & layer_0[11038]); 
    assign out[5065] = layer_0[1058] ^ layer_0[10417]; 
    assign out[5066] = layer_0[817] ^ layer_0[7122]; 
    assign out[5067] = ~(layer_0[8880] ^ layer_0[7401]); 
    assign out[5068] = ~(layer_0[6888] ^ layer_0[102]); 
    assign out[5069] = layer_0[11399]; 
    assign out[5070] = layer_0[11106] ^ layer_0[3935]; 
    assign out[5071] = layer_0[272] ^ layer_0[1267]; 
    assign out[5072] = layer_0[3441]; 
    assign out[5073] = ~(layer_0[9855] ^ layer_0[5482]); 
    assign out[5074] = layer_0[144] ^ layer_0[1469]; 
    assign out[5075] = ~(layer_0[4150] ^ layer_0[8513]); 
    assign out[5076] = layer_0[3261] ^ layer_0[2719]; 
    assign out[5077] = layer_0[5984] ^ layer_0[3414]; 
    assign out[5078] = ~(layer_0[4403] & layer_0[652]); 
    assign out[5079] = ~layer_0[3192] | (layer_0[8101] & layer_0[3192]); 
    assign out[5080] = layer_0[5554] ^ layer_0[4877]; 
    assign out[5081] = layer_0[4471] ^ layer_0[5022]; 
    assign out[5082] = ~layer_0[9293] | (layer_0[9293] & layer_0[2722]); 
    assign out[5083] = layer_0[9292]; 
    assign out[5084] = layer_0[7559] ^ layer_0[11096]; 
    assign out[5085] = ~layer_0[7383]; 
    assign out[5086] = layer_0[8879]; 
    assign out[5087] = layer_0[11179] ^ layer_0[5106]; 
    assign out[5088] = ~layer_0[9012]; 
    assign out[5089] = ~layer_0[2993]; 
    assign out[5090] = layer_0[1887] ^ layer_0[7215]; 
    assign out[5091] = ~(layer_0[1000] ^ layer_0[9705]); 
    assign out[5092] = ~layer_0[2470]; 
    assign out[5093] = ~(layer_0[8833] ^ layer_0[5487]); 
    assign out[5094] = layer_0[8059] & ~layer_0[8084]; 
    assign out[5095] = ~(layer_0[11673] ^ layer_0[2010]); 
    assign out[5096] = layer_0[11377] & layer_0[11068]; 
    assign out[5097] = layer_0[5230] | layer_0[4880]; 
    assign out[5098] = ~(layer_0[7534] ^ layer_0[7661]); 
    assign out[5099] = ~(layer_0[5333] ^ layer_0[5207]); 
    assign out[5100] = ~(layer_0[4322] ^ layer_0[10421]); 
    assign out[5101] = ~layer_0[9700]; 
    assign out[5102] = layer_0[391] ^ layer_0[4834]; 
    assign out[5103] = layer_0[107] ^ layer_0[6380]; 
    assign out[5104] = ~layer_0[3616]; 
    assign out[5105] = layer_0[6879]; 
    assign out[5106] = layer_0[2657] ^ layer_0[9875]; 
    assign out[5107] = ~(layer_0[10101] ^ layer_0[11986]); 
    assign out[5108] = layer_0[3030]; 
    assign out[5109] = layer_0[10912]; 
    assign out[5110] = ~layer_0[1529]; 
    assign out[5111] = layer_0[11395] | layer_0[3024]; 
    assign out[5112] = layer_0[3227]; 
    assign out[5113] = ~layer_0[2873] | (layer_0[9479] & layer_0[2873]); 
    assign out[5114] = ~(layer_0[6276] ^ layer_0[6603]); 
    assign out[5115] = layer_0[4704] & ~layer_0[8708]; 
    assign out[5116] = ~(layer_0[10719] | layer_0[3156]); 
    assign out[5117] = layer_0[9513]; 
    assign out[5118] = ~(layer_0[1701] ^ layer_0[11730]); 
    assign out[5119] = ~layer_0[8927]; 
    assign out[5120] = ~(layer_0[9635] ^ layer_0[390]); 
    assign out[5121] = ~layer_0[2097]; 
    assign out[5122] = ~(layer_0[1029] ^ layer_0[173]); 
    assign out[5123] = layer_0[2684] ^ layer_0[7389]; 
    assign out[5124] = ~layer_0[3066]; 
    assign out[5125] = ~(layer_0[8145] & layer_0[378]); 
    assign out[5126] = ~layer_0[1209] | (layer_0[1363] & layer_0[1209]); 
    assign out[5127] = ~(layer_0[3178] ^ layer_0[5536]); 
    assign out[5128] = ~layer_0[3184]; 
    assign out[5129] = ~(layer_0[1702] ^ layer_0[11229]); 
    assign out[5130] = layer_0[8077] ^ layer_0[5582]; 
    assign out[5131] = layer_0[11187] ^ layer_0[740]; 
    assign out[5132] = layer_0[7495] ^ layer_0[3639]; 
    assign out[5133] = ~(layer_0[8467] ^ layer_0[893]); 
    assign out[5134] = layer_0[1013] & ~layer_0[3022]; 
    assign out[5135] = ~layer_0[3789]; 
    assign out[5136] = ~(layer_0[232] ^ layer_0[8815]); 
    assign out[5137] = ~(layer_0[9149] | layer_0[1390]); 
    assign out[5138] = layer_0[6356] ^ layer_0[1285]; 
    assign out[5139] = layer_0[5192] ^ layer_0[9248]; 
    assign out[5140] = ~layer_0[8241] | (layer_0[8241] & layer_0[11745]); 
    assign out[5141] = layer_0[11625] & layer_0[6559]; 
    assign out[5142] = ~(layer_0[8840] ^ layer_0[4132]); 
    assign out[5143] = layer_0[10059] ^ layer_0[288]; 
    assign out[5144] = ~(layer_0[206] ^ layer_0[4582]); 
    assign out[5145] = layer_0[5125] ^ layer_0[6897]; 
    assign out[5146] = ~(layer_0[6158] ^ layer_0[3132]); 
    assign out[5147] = layer_0[7754] ^ layer_0[1978]; 
    assign out[5148] = layer_0[11330] ^ layer_0[6435]; 
    assign out[5149] = layer_0[11188] ^ layer_0[5234]; 
    assign out[5150] = ~(layer_0[3730] ^ layer_0[10709]); 
    assign out[5151] = ~(layer_0[6918] ^ layer_0[2437]); 
    assign out[5152] = layer_0[2077] ^ layer_0[9725]; 
    assign out[5153] = layer_0[10825]; 
    assign out[5154] = layer_0[5444] ^ layer_0[8102]; 
    assign out[5155] = layer_0[9970] ^ layer_0[4735]; 
    assign out[5156] = ~(layer_0[4932] ^ layer_0[7371]); 
    assign out[5157] = ~(layer_0[6770] & layer_0[281]); 
    assign out[5158] = layer_0[6000] ^ layer_0[2883]; 
    assign out[5159] = layer_0[381] ^ layer_0[4379]; 
    assign out[5160] = ~(layer_0[5912] & layer_0[10732]); 
    assign out[5161] = layer_0[732] ^ layer_0[7731]; 
    assign out[5162] = layer_0[99]; 
    assign out[5163] = layer_0[5669] & ~layer_0[7370]; 
    assign out[5164] = ~layer_0[1112]; 
    assign out[5165] = layer_0[1433] ^ layer_0[4338]; 
    assign out[5166] = ~(layer_0[11657] ^ layer_0[1294]); 
    assign out[5167] = layer_0[8365] ^ layer_0[4504]; 
    assign out[5168] = layer_0[629] ^ layer_0[5216]; 
    assign out[5169] = layer_0[3548] | layer_0[3598]; 
    assign out[5170] = layer_0[9820] ^ layer_0[7723]; 
    assign out[5171] = layer_0[5775] & ~layer_0[5949]; 
    assign out[5172] = layer_0[6799] ^ layer_0[472]; 
    assign out[5173] = ~(layer_0[5028] & layer_0[3821]); 
    assign out[5174] = ~(layer_0[3871] ^ layer_0[2186]); 
    assign out[5175] = layer_0[770] & ~layer_0[1446]; 
    assign out[5176] = layer_0[2414] & ~layer_0[8041]; 
    assign out[5177] = layer_0[10083]; 
    assign out[5178] = layer_0[9379] ^ layer_0[10219]; 
    assign out[5179] = ~(layer_0[7591] ^ layer_0[1927]); 
    assign out[5180] = ~(layer_0[5820] ^ layer_0[3928]); 
    assign out[5181] = ~(layer_0[9245] ^ layer_0[1896]); 
    assign out[5182] = ~(layer_0[678] ^ layer_0[11737]); 
    assign out[5183] = layer_0[4031] ^ layer_0[4656]; 
    assign out[5184] = ~layer_0[9495] | (layer_0[1199] & layer_0[9495]); 
    assign out[5185] = layer_0[867] & layer_0[6491]; 
    assign out[5186] = ~(layer_0[3718] ^ layer_0[10245]); 
    assign out[5187] = ~(layer_0[7913] ^ layer_0[2688]); 
    assign out[5188] = ~(layer_0[11174] ^ layer_0[4681]); 
    assign out[5189] = layer_0[1015] & ~layer_0[10420]; 
    assign out[5190] = layer_0[6081] ^ layer_0[2690]; 
    assign out[5191] = ~layer_0[8093] | (layer_0[8093] & layer_0[2666]); 
    assign out[5192] = layer_0[6484] ^ layer_0[11735]; 
    assign out[5193] = layer_0[8164]; 
    assign out[5194] = ~layer_0[11175] | (layer_0[11175] & layer_0[9937]); 
    assign out[5195] = layer_0[6422] ^ layer_0[3602]; 
    assign out[5196] = layer_0[155] & ~layer_0[4550]; 
    assign out[5197] = layer_0[1289] & ~layer_0[1380]; 
    assign out[5198] = ~(layer_0[9045] ^ layer_0[2992]); 
    assign out[5199] = layer_0[2151] & ~layer_0[6893]; 
    assign out[5200] = layer_0[2170]; 
    assign out[5201] = ~layer_0[3201] | (layer_0[6719] & layer_0[3201]); 
    assign out[5202] = layer_0[5872] ^ layer_0[1076]; 
    assign out[5203] = ~layer_0[8761]; 
    assign out[5204] = layer_0[6091] ^ layer_0[955]; 
    assign out[5205] = ~(layer_0[8491] ^ layer_0[2798]); 
    assign out[5206] = layer_0[9783] ^ layer_0[6846]; 
    assign out[5207] = layer_0[1613] & layer_0[1070]; 
    assign out[5208] = layer_0[1079] ^ layer_0[9202]; 
    assign out[5209] = ~(layer_0[10534] ^ layer_0[924]); 
    assign out[5210] = ~(layer_0[5231] ^ layer_0[7647]); 
    assign out[5211] = layer_0[5052] ^ layer_0[3384]; 
    assign out[5212] = layer_0[5481] & ~layer_0[928]; 
    assign out[5213] = ~(layer_0[794] ^ layer_0[533]); 
    assign out[5214] = ~layer_0[3657] | (layer_0[1852] & layer_0[3657]); 
    assign out[5215] = layer_0[4869] ^ layer_0[5641]; 
    assign out[5216] = layer_0[2852] ^ layer_0[11102]; 
    assign out[5217] = ~layer_0[6922]; 
    assign out[5218] = ~(layer_0[2987] ^ layer_0[8803]); 
    assign out[5219] = layer_0[7506] ^ layer_0[8821]; 
    assign out[5220] = ~(layer_0[3600] & layer_0[307]); 
    assign out[5221] = layer_0[9222]; 
    assign out[5222] = layer_0[6727] ^ layer_0[7161]; 
    assign out[5223] = ~(layer_0[4498] & layer_0[2704]); 
    assign out[5224] = ~(layer_0[896] ^ layer_0[1325]); 
    assign out[5225] = layer_0[8070] ^ layer_0[6323]; 
    assign out[5226] = layer_0[4222] ^ layer_0[10542]; 
    assign out[5227] = ~layer_0[3936]; 
    assign out[5228] = ~(layer_0[11250] ^ layer_0[8788]); 
    assign out[5229] = layer_0[6654] ^ layer_0[8598]; 
    assign out[5230] = layer_0[4827] | layer_0[1544]; 
    assign out[5231] = ~layer_0[3154]; 
    assign out[5232] = ~(layer_0[7205] ^ layer_0[1262]); 
    assign out[5233] = ~(layer_0[3260] ^ layer_0[10323]); 
    assign out[5234] = ~(layer_0[4182] | layer_0[8863]); 
    assign out[5235] = ~(layer_0[4878] & layer_0[8481]); 
    assign out[5236] = ~(layer_0[6655] ^ layer_0[2830]); 
    assign out[5237] = ~(layer_0[1913] ^ layer_0[11140]); 
    assign out[5238] = layer_0[6826] ^ layer_0[10940]; 
    assign out[5239] = ~(layer_0[10823] ^ layer_0[10831]); 
    assign out[5240] = ~layer_0[10224]; 
    assign out[5241] = ~(layer_0[10512] | layer_0[4115]); 
    assign out[5242] = ~layer_0[10344]; 
    assign out[5243] = ~(layer_0[6245] ^ layer_0[9612]); 
    assign out[5244] = ~layer_0[3246]; 
    assign out[5245] = ~layer_0[8045] | (layer_0[8045] & layer_0[9997]); 
    assign out[5246] = ~layer_0[2938] | (layer_0[2938] & layer_0[9267]); 
    assign out[5247] = ~(layer_0[3610] ^ layer_0[1838]); 
    assign out[5248] = layer_0[7960] ^ layer_0[2603]; 
    assign out[5249] = layer_0[8102] ^ layer_0[930]; 
    assign out[5250] = ~layer_0[3329] | (layer_0[3329] & layer_0[11752]); 
    assign out[5251] = ~(layer_0[10865] ^ layer_0[10934]); 
    assign out[5252] = layer_0[2686] ^ layer_0[2356]; 
    assign out[5253] = ~layer_0[9360]; 
    assign out[5254] = layer_0[11201] | layer_0[5972]; 
    assign out[5255] = layer_0[7449] ^ layer_0[10851]; 
    assign out[5256] = ~(layer_0[1052] & layer_0[4729]); 
    assign out[5257] = layer_0[5449] | layer_0[676]; 
    assign out[5258] = layer_0[7194] & ~layer_0[7973]; 
    assign out[5259] = ~(layer_0[6583] ^ layer_0[7726]); 
    assign out[5260] = ~(layer_0[630] ^ layer_0[476]); 
    assign out[5261] = ~(layer_0[6596] ^ layer_0[2780]); 
    assign out[5262] = layer_0[1073]; 
    assign out[5263] = ~(layer_0[8891] & layer_0[7961]); 
    assign out[5264] = ~layer_0[11263] | (layer_0[2595] & layer_0[11263]); 
    assign out[5265] = layer_0[3902] ^ layer_0[458]; 
    assign out[5266] = layer_0[8629] ^ layer_0[8392]; 
    assign out[5267] = ~(layer_0[5948] ^ layer_0[8754]); 
    assign out[5268] = ~layer_0[10167] | (layer_0[10167] & layer_0[2648]); 
    assign out[5269] = ~(layer_0[4699] ^ layer_0[7543]); 
    assign out[5270] = layer_0[3721]; 
    assign out[5271] = layer_0[8936] & ~layer_0[10577]; 
    assign out[5272] = layer_0[4251]; 
    assign out[5273] = ~(layer_0[1352] ^ layer_0[3961]); 
    assign out[5274] = layer_0[1930] | layer_0[6142]; 
    assign out[5275] = ~layer_0[5852] | (layer_0[2786] & layer_0[5852]); 
    assign out[5276] = layer_0[6804]; 
    assign out[5277] = ~layer_0[10927] | (layer_0[8273] & layer_0[10927]); 
    assign out[5278] = ~(layer_0[10798] ^ layer_0[11934]); 
    assign out[5279] = layer_0[3476] ^ layer_0[5484]; 
    assign out[5280] = ~(layer_0[1636] ^ layer_0[7571]); 
    assign out[5281] = layer_0[11248] & layer_0[2485]; 
    assign out[5282] = ~layer_0[6239]; 
    assign out[5283] = layer_0[9567] & ~layer_0[10123]; 
    assign out[5284] = ~(layer_0[10303] ^ layer_0[9898]); 
    assign out[5285] = layer_0[8555] ^ layer_0[11541]; 
    assign out[5286] = layer_0[6138] ^ layer_0[8414]; 
    assign out[5287] = ~(layer_0[5563] ^ layer_0[11940]); 
    assign out[5288] = layer_0[7359] & ~layer_0[752]; 
    assign out[5289] = layer_0[7314] & ~layer_0[7715]; 
    assign out[5290] = ~(layer_0[5040] & layer_0[9129]); 
    assign out[5291] = ~(layer_0[10565] ^ layer_0[5316]); 
    assign out[5292] = ~(layer_0[6088] ^ layer_0[8862]); 
    assign out[5293] = layer_0[3977] ^ layer_0[5760]; 
    assign out[5294] = ~layer_0[5322]; 
    assign out[5295] = layer_0[8566] ^ layer_0[6809]; 
    assign out[5296] = layer_0[2782] ^ layer_0[10937]; 
    assign out[5297] = ~(layer_0[5568] ^ layer_0[9880]); 
    assign out[5298] = layer_0[9411] ^ layer_0[4542]; 
    assign out[5299] = ~(layer_0[3411] & layer_0[3139]); 
    assign out[5300] = ~(layer_0[4414] ^ layer_0[11399]); 
    assign out[5301] = ~(layer_0[9076] ^ layer_0[11732]); 
    assign out[5302] = ~(layer_0[4372] & layer_0[8463]); 
    assign out[5303] = ~(layer_0[10401] ^ layer_0[11460]); 
    assign out[5304] = layer_0[6857] | layer_0[10467]; 
    assign out[5305] = layer_0[11838] & ~layer_0[1517]; 
    assign out[5306] = ~(layer_0[6018] ^ layer_0[1831]); 
    assign out[5307] = ~(layer_0[2436] ^ layer_0[1027]); 
    assign out[5308] = ~(layer_0[11614] ^ layer_0[6062]); 
    assign out[5309] = layer_0[6894] ^ layer_0[1508]; 
    assign out[5310] = ~layer_0[3495]; 
    assign out[5311] = layer_0[1663]; 
    assign out[5312] = ~layer_0[8799] | (layer_0[8799] & layer_0[4659]); 
    assign out[5313] = layer_0[7900] & layer_0[9944]; 
    assign out[5314] = layer_0[1276] ^ layer_0[4298]; 
    assign out[5315] = layer_0[7217] ^ layer_0[1001]; 
    assign out[5316] = ~layer_0[712]; 
    assign out[5317] = layer_0[10748] ^ layer_0[8926]; 
    assign out[5318] = ~(layer_0[215] ^ layer_0[899]); 
    assign out[5319] = layer_0[8030] | layer_0[5626]; 
    assign out[5320] = layer_0[6534] ^ layer_0[2312]; 
    assign out[5321] = layer_0[8989] & ~layer_0[622]; 
    assign out[5322] = ~layer_0[4172]; 
    assign out[5323] = ~(layer_0[5190] ^ layer_0[9680]); 
    assign out[5324] = ~layer_0[332]; 
    assign out[5325] = layer_0[4030] | layer_0[10288]; 
    assign out[5326] = layer_0[5105] ^ layer_0[9840]; 
    assign out[5327] = layer_0[11500] & ~layer_0[7606]; 
    assign out[5328] = layer_0[6371] ^ layer_0[5263]; 
    assign out[5329] = layer_0[6882] & ~layer_0[854]; 
    assign out[5330] = layer_0[2818]; 
    assign out[5331] = layer_0[7113] ^ layer_0[1960]; 
    assign out[5332] = ~(layer_0[4953] ^ layer_0[967]); 
    assign out[5333] = ~layer_0[5529]; 
    assign out[5334] = ~(layer_0[192] ^ layer_0[7477]); 
    assign out[5335] = ~(layer_0[753] ^ layer_0[7942]); 
    assign out[5336] = layer_0[66] ^ layer_0[2371]; 
    assign out[5337] = layer_0[11287] ^ layer_0[6867]; 
    assign out[5338] = ~layer_0[8313] | (layer_0[8313] & layer_0[8034]); 
    assign out[5339] = ~(layer_0[1069] ^ layer_0[8037]); 
    assign out[5340] = layer_0[5016] ^ layer_0[2318]; 
    assign out[5341] = ~(layer_0[5309] ^ layer_0[4276]); 
    assign out[5342] = ~(layer_0[1277] ^ layer_0[7114]); 
    assign out[5343] = ~layer_0[7604]; 
    assign out[5344] = ~(layer_0[7797] | layer_0[5845]); 
    assign out[5345] = ~layer_0[9023]; 
    assign out[5346] = layer_0[8619] ^ layer_0[5491]; 
    assign out[5347] = ~(layer_0[8184] ^ layer_0[8261]); 
    assign out[5348] = ~layer_0[800]; 
    assign out[5349] = layer_0[2687] ^ layer_0[3409]; 
    assign out[5350] = layer_0[7190] | layer_0[6408]; 
    assign out[5351] = ~(layer_0[7629] | layer_0[9425]); 
    assign out[5352] = layer_0[612]; 
    assign out[5353] = ~(layer_0[10839] & layer_0[8526]); 
    assign out[5354] = ~(layer_0[1790] ^ layer_0[5206]); 
    assign out[5355] = layer_0[2311] & ~layer_0[3297]; 
    assign out[5356] = layer_0[2218] ^ layer_0[10863]; 
    assign out[5357] = ~(layer_0[2609] ^ layer_0[11618]); 
    assign out[5358] = layer_0[2095] ^ layer_0[6529]; 
    assign out[5359] = layer_0[9665] ^ layer_0[5962]; 
    assign out[5360] = ~(layer_0[2751] ^ layer_0[8771]); 
    assign out[5361] = ~layer_0[11367]; 
    assign out[5362] = ~(layer_0[8353] ^ layer_0[5088]); 
    assign out[5363] = ~layer_0[11317] | (layer_0[11317] & layer_0[8910]); 
    assign out[5364] = layer_0[9484] ^ layer_0[11917]; 
    assign out[5365] = layer_0[8836] ^ layer_0[11532]; 
    assign out[5366] = layer_0[11999] ^ layer_0[11114]; 
    assign out[5367] = layer_0[7709] ^ layer_0[3599]; 
    assign out[5368] = ~(layer_0[5298] ^ layer_0[4561]); 
    assign out[5369] = layer_0[7645]; 
    assign out[5370] = layer_0[1947] ^ layer_0[11293]; 
    assign out[5371] = layer_0[1724] ^ layer_0[11369]; 
    assign out[5372] = layer_0[1189]; 
    assign out[5373] = layer_0[10943] ^ layer_0[4862]; 
    assign out[5374] = ~(layer_0[4569] ^ layer_0[3676]); 
    assign out[5375] = ~(layer_0[11301] | layer_0[1681]); 
    assign out[5376] = ~(layer_0[5076] ^ layer_0[10538]); 
    assign out[5377] = layer_0[4497] ^ layer_0[9941]; 
    assign out[5378] = ~layer_0[3795] | (layer_0[6853] & layer_0[3795]); 
    assign out[5379] = ~(layer_0[7236] ^ layer_0[6802]); 
    assign out[5380] = ~(layer_0[5308] ^ layer_0[6318]); 
    assign out[5381] = layer_0[9518] ^ layer_0[882]; 
    assign out[5382] = layer_0[36] & ~layer_0[9667]; 
    assign out[5383] = layer_0[1967] | layer_0[8757]; 
    assign out[5384] = layer_0[8464] ^ layer_0[9113]; 
    assign out[5385] = layer_0[9258] ^ layer_0[11814]; 
    assign out[5386] = layer_0[7750] ^ layer_0[8517]; 
    assign out[5387] = layer_0[6052] & ~layer_0[10271]; 
    assign out[5388] = ~layer_0[1459] | (layer_0[8661] & layer_0[1459]); 
    assign out[5389] = layer_0[10791] ^ layer_0[2105]; 
    assign out[5390] = ~layer_0[6161]; 
    assign out[5391] = layer_0[9278] ^ layer_0[9877]; 
    assign out[5392] = layer_0[319]; 
    assign out[5393] = ~(layer_0[540] ^ layer_0[2416]); 
    assign out[5394] = layer_0[11274] ^ layer_0[1252]; 
    assign out[5395] = ~(layer_0[865] ^ layer_0[11049]); 
    assign out[5396] = ~(layer_0[7749] ^ layer_0[9771]); 
    assign out[5397] = layer_0[6131] & layer_0[3692]; 
    assign out[5398] = layer_0[6146]; 
    assign out[5399] = layer_0[900] ^ layer_0[895]; 
    assign out[5400] = ~(layer_0[11319] | layer_0[10869]); 
    assign out[5401] = layer_0[6051] ^ layer_0[3508]; 
    assign out[5402] = layer_0[4823] ^ layer_0[8673]; 
    assign out[5403] = ~layer_0[2404]; 
    assign out[5404] = ~layer_0[10472]; 
    assign out[5405] = ~(layer_0[448] & layer_0[6689]); 
    assign out[5406] = ~(layer_0[3841] | layer_0[29]); 
    assign out[5407] = layer_0[10498] ^ layer_0[11449]; 
    assign out[5408] = layer_0[7630] | layer_0[2728]; 
    assign out[5409] = layer_0[5398] ^ layer_0[11581]; 
    assign out[5410] = ~layer_0[6625]; 
    assign out[5411] = ~(layer_0[8645] ^ layer_0[2516]); 
    assign out[5412] = layer_0[7638] & ~layer_0[11390]; 
    assign out[5413] = ~(layer_0[11602] ^ layer_0[5131]); 
    assign out[5414] = ~layer_0[3680] | (layer_0[8779] & layer_0[3680]); 
    assign out[5415] = ~(layer_0[105] ^ layer_0[7743]); 
    assign out[5416] = layer_0[10341] & layer_0[5586]; 
    assign out[5417] = ~(layer_0[10539] ^ layer_0[11144]); 
    assign out[5418] = layer_0[5042]; 
    assign out[5419] = ~(layer_0[1733] ^ layer_0[9192]); 
    assign out[5420] = layer_0[6992] ^ layer_0[274]; 
    assign out[5421] = ~layer_0[10931] | (layer_0[10931] & layer_0[7538]); 
    assign out[5422] = ~layer_0[10427]; 
    assign out[5423] = layer_0[2021] ^ layer_0[3824]; 
    assign out[5424] = layer_0[6187]; 
    assign out[5425] = ~layer_0[11338]; 
    assign out[5426] = ~(layer_0[11622] ^ layer_0[11124]); 
    assign out[5427] = ~layer_0[11697] | (layer_0[11697] & layer_0[309]); 
    assign out[5428] = layer_0[5607] ^ layer_0[6292]; 
    assign out[5429] = layer_0[9404] ^ layer_0[8857]; 
    assign out[5430] = layer_0[11991]; 
    assign out[5431] = layer_0[8668] | layer_0[75]; 
    assign out[5432] = layer_0[11986] & ~layer_0[1082]; 
    assign out[5433] = layer_0[8686] ^ layer_0[1119]; 
    assign out[5434] = layer_0[6935] ^ layer_0[8918]; 
    assign out[5435] = layer_0[4421]; 
    assign out[5436] = layer_0[86] ^ layer_0[8910]; 
    assign out[5437] = layer_0[507] ^ layer_0[6362]; 
    assign out[5438] = layer_0[7027] & ~layer_0[4044]; 
    assign out[5439] = ~layer_0[6034]; 
    assign out[5440] = ~(layer_0[6122] | layer_0[7684]); 
    assign out[5441] = layer_0[9584] ^ layer_0[8190]; 
    assign out[5442] = ~layer_0[800]; 
    assign out[5443] = layer_0[11972]; 
    assign out[5444] = layer_0[1301] ^ layer_0[4507]; 
    assign out[5445] = layer_0[9473] ^ layer_0[11203]; 
    assign out[5446] = layer_0[1147] & layer_0[9328]; 
    assign out[5447] = ~(layer_0[890] ^ layer_0[4086]); 
    assign out[5448] = layer_0[4604] ^ layer_0[2239]; 
    assign out[5449] = layer_0[10717] ^ layer_0[6842]; 
    assign out[5450] = layer_0[2023]; 
    assign out[5451] = layer_0[11769]; 
    assign out[5452] = layer_0[1478] ^ layer_0[2904]; 
    assign out[5453] = ~(layer_0[8169] ^ layer_0[4311]); 
    assign out[5454] = ~layer_0[11688] | (layer_0[3987] & layer_0[11688]); 
    assign out[5455] = layer_0[11268] | layer_0[10622]; 
    assign out[5456] = layer_0[2389] & ~layer_0[3401]; 
    assign out[5457] = ~(layer_0[11669] ^ layer_0[231]); 
    assign out[5458] = layer_0[11017] ^ layer_0[9045]; 
    assign out[5459] = ~layer_0[6925]; 
    assign out[5460] = ~(layer_0[5563] ^ layer_0[10982]); 
    assign out[5461] = ~(layer_0[11713] ^ layer_0[10138]); 
    assign out[5462] = ~layer_0[11775]; 
    assign out[5463] = ~(layer_0[3189] & layer_0[6093]); 
    assign out[5464] = ~layer_0[3182]; 
    assign out[5465] = ~(layer_0[11591] ^ layer_0[4596]); 
    assign out[5466] = ~layer_0[4925]; 
    assign out[5467] = ~(layer_0[9650] ^ layer_0[6976]); 
    assign out[5468] = layer_0[11699] & layer_0[9154]; 
    assign out[5469] = layer_0[4840]; 
    assign out[5470] = ~layer_0[2133]; 
    assign out[5471] = ~(layer_0[1641] ^ layer_0[842]); 
    assign out[5472] = layer_0[11138] ^ layer_0[11487]; 
    assign out[5473] = ~(layer_0[255] ^ layer_0[10944]); 
    assign out[5474] = ~(layer_0[11924] & layer_0[644]); 
    assign out[5475] = layer_0[11512] ^ layer_0[6865]; 
    assign out[5476] = layer_0[2806] ^ layer_0[4696]; 
    assign out[5477] = layer_0[636] ^ layer_0[3276]; 
    assign out[5478] = ~layer_0[2843] | (layer_0[2843] & layer_0[533]); 
    assign out[5479] = ~(layer_0[10572] ^ layer_0[6805]); 
    assign out[5480] = ~(layer_0[9390] ^ layer_0[2620]); 
    assign out[5481] = ~(layer_0[10085] ^ layer_0[5193]); 
    assign out[5482] = layer_0[586] ^ layer_0[2297]; 
    assign out[5483] = layer_0[3776] ^ layer_0[939]; 
    assign out[5484] = layer_0[10717] | layer_0[4014]; 
    assign out[5485] = ~(layer_0[4970] & layer_0[10761]); 
    assign out[5486] = layer_0[10364] & layer_0[4676]; 
    assign out[5487] = ~(layer_0[2257] | layer_0[6707]); 
    assign out[5488] = ~(layer_0[7983] ^ layer_0[4371]); 
    assign out[5489] = layer_0[2185] ^ layer_0[11093]; 
    assign out[5490] = ~(layer_0[9203] ^ layer_0[3307]); 
    assign out[5491] = ~(layer_0[1130] ^ layer_0[3050]); 
    assign out[5492] = layer_0[9952]; 
    assign out[5493] = ~(layer_0[10480] | layer_0[6301]); 
    assign out[5494] = ~(layer_0[4657] & layer_0[2594]); 
    assign out[5495] = layer_0[3095] | layer_0[5940]; 
    assign out[5496] = layer_0[3570] ^ layer_0[1673]; 
    assign out[5497] = ~(layer_0[2995] ^ layer_0[1982]); 
    assign out[5498] = layer_0[5144] ^ layer_0[181]; 
    assign out[5499] = ~(layer_0[3828] ^ layer_0[4215]); 
    assign out[5500] = layer_0[983] & ~layer_0[7954]; 
    assign out[5501] = layer_0[7184] ^ layer_0[7569]; 
    assign out[5502] = ~(layer_0[11756] ^ layer_0[9704]); 
    assign out[5503] = ~(layer_0[6206] ^ layer_0[6943]); 
    assign out[5504] = layer_0[9562] | layer_0[7798]; 
    assign out[5505] = ~layer_0[955] | (layer_0[3898] & layer_0[955]); 
    assign out[5506] = layer_0[9602] & ~layer_0[4171]; 
    assign out[5507] = ~layer_0[9175]; 
    assign out[5508] = ~(layer_0[9248] ^ layer_0[6024]); 
    assign out[5509] = ~(layer_0[5332] ^ layer_0[3751]); 
    assign out[5510] = ~(layer_0[1837] ^ layer_0[6896]); 
    assign out[5511] = layer_0[1395]; 
    assign out[5512] = ~(layer_0[6576] ^ layer_0[11874]); 
    assign out[5513] = ~(layer_0[9989] ^ layer_0[5647]); 
    assign out[5514] = ~layer_0[1683] | (layer_0[9972] & layer_0[1683]); 
    assign out[5515] = ~(layer_0[5710] ^ layer_0[11261]); 
    assign out[5516] = ~layer_0[5986]; 
    assign out[5517] = layer_0[11973] ^ layer_0[366]; 
    assign out[5518] = ~(layer_0[10416] ^ layer_0[11611]); 
    assign out[5519] = layer_0[4891] ^ layer_0[9079]; 
    assign out[5520] = layer_0[9059] ^ layer_0[648]; 
    assign out[5521] = ~layer_0[11777] | (layer_0[3589] & layer_0[11777]); 
    assign out[5522] = layer_0[7254] ^ layer_0[4052]; 
    assign out[5523] = ~(layer_0[3404] | layer_0[10808]); 
    assign out[5524] = ~layer_0[5455]; 
    assign out[5525] = layer_0[8837] ^ layer_0[9601]; 
    assign out[5526] = layer_0[8340] ^ layer_0[6012]; 
    assign out[5527] = ~(layer_0[9849] ^ layer_0[10879]); 
    assign out[5528] = layer_0[1024] ^ layer_0[11447]; 
    assign out[5529] = ~(layer_0[3394] ^ layer_0[3712]); 
    assign out[5530] = ~(layer_0[5749] ^ layer_0[11423]); 
    assign out[5531] = layer_0[11619] ^ layer_0[1688]; 
    assign out[5532] = ~(layer_0[942] ^ layer_0[7251]); 
    assign out[5533] = ~layer_0[445]; 
    assign out[5534] = layer_0[3622] ^ layer_0[8393]; 
    assign out[5535] = ~(layer_0[5082] ^ layer_0[5277]); 
    assign out[5536] = ~(layer_0[4483] ^ layer_0[6021]); 
    assign out[5537] = ~(layer_0[9804] ^ layer_0[544]); 
    assign out[5538] = layer_0[8762] ^ layer_0[10941]; 
    assign out[5539] = layer_0[407] ^ layer_0[7345]; 
    assign out[5540] = ~(layer_0[4422] ^ layer_0[11009]); 
    assign out[5541] = layer_0[5847]; 
    assign out[5542] = ~(layer_0[6754] ^ layer_0[9587]); 
    assign out[5543] = layer_0[8746] ^ layer_0[11018]; 
    assign out[5544] = layer_0[11053] ^ layer_0[9431]; 
    assign out[5545] = layer_0[9712] & ~layer_0[7433]; 
    assign out[5546] = ~(layer_0[6199] ^ layer_0[4342]); 
    assign out[5547] = ~(layer_0[2755] ^ layer_0[6519]); 
    assign out[5548] = layer_0[9472] & layer_0[9063]; 
    assign out[5549] = layer_0[7796]; 
    assign out[5550] = layer_0[2229] ^ layer_0[4219]; 
    assign out[5551] = ~(layer_0[2311] ^ layer_0[9466]); 
    assign out[5552] = ~(layer_0[5908] ^ layer_0[5615]); 
    assign out[5553] = layer_0[1299] ^ layer_0[1369]; 
    assign out[5554] = ~(layer_0[11042] ^ layer_0[8425]); 
    assign out[5555] = layer_0[4162] & ~layer_0[6687]; 
    assign out[5556] = ~(layer_0[4487] & layer_0[11922]); 
    assign out[5557] = ~layer_0[6155]; 
    assign out[5558] = layer_0[3989]; 
    assign out[5559] = ~(layer_0[9388] ^ layer_0[8140]); 
    assign out[5560] = ~(layer_0[4451] ^ layer_0[5705]); 
    assign out[5561] = ~layer_0[8993] | (layer_0[8993] & layer_0[3930]); 
    assign out[5562] = ~layer_0[92] | (layer_0[6354] & layer_0[92]); 
    assign out[5563] = ~(layer_0[5179] & layer_0[11169]); 
    assign out[5564] = layer_0[2964] ^ layer_0[10155]; 
    assign out[5565] = ~(layer_0[9386] ^ layer_0[8062]); 
    assign out[5566] = ~layer_0[8987] | (layer_0[8987] & layer_0[1497]); 
    assign out[5567] = ~(layer_0[6570] & layer_0[5866]); 
    assign out[5568] = layer_0[4617]; 
    assign out[5569] = layer_0[434] ^ layer_0[11898]; 
    assign out[5570] = ~(layer_0[10783] ^ layer_0[4746]); 
    assign out[5571] = ~(layer_0[5794] | layer_0[9367]); 
    assign out[5572] = ~layer_0[3748]; 
    assign out[5573] = ~(layer_0[2427] ^ layer_0[10749]); 
    assign out[5574] = layer_0[7309] ^ layer_0[9209]; 
    assign out[5575] = layer_0[6290]; 
    assign out[5576] = layer_0[11310] ^ layer_0[2206]; 
    assign out[5577] = ~(layer_0[2132] | layer_0[6982]); 
    assign out[5578] = ~(layer_0[2605] ^ layer_0[934]); 
    assign out[5579] = ~(layer_0[11876] ^ layer_0[9979]); 
    assign out[5580] = ~layer_0[985]; 
    assign out[5581] = layer_0[3788] ^ layer_0[1288]; 
    assign out[5582] = ~(layer_0[7177] ^ layer_0[2705]); 
    assign out[5583] = ~(layer_0[9375] ^ layer_0[9474]); 
    assign out[5584] = ~layer_0[1224]; 
    assign out[5585] = layer_0[6676] ^ layer_0[3513]; 
    assign out[5586] = layer_0[9627] ^ layer_0[2903]; 
    assign out[5587] = ~(layer_0[3596] & layer_0[6074]); 
    assign out[5588] = layer_0[3832] ^ layer_0[11680]; 
    assign out[5589] = ~(layer_0[9253] ^ layer_0[5013]); 
    assign out[5590] = ~layer_0[6613]; 
    assign out[5591] = ~(layer_0[3287] | layer_0[7407]); 
    assign out[5592] = ~(layer_0[1173] ^ layer_0[10631]); 
    assign out[5593] = ~(layer_0[1084] ^ layer_0[10218]); 
    assign out[5594] = ~(layer_0[5555] ^ layer_0[440]); 
    assign out[5595] = layer_0[8693] ^ layer_0[9917]; 
    assign out[5596] = layer_0[1575] ^ layer_0[6661]; 
    assign out[5597] = layer_0[6468] & ~layer_0[10301]; 
    assign out[5598] = ~layer_0[5084]; 
    assign out[5599] = layer_0[7634]; 
    assign out[5600] = ~(layer_0[8876] ^ layer_0[6190]); 
    assign out[5601] = ~(layer_0[7701] ^ layer_0[2343]); 
    assign out[5602] = ~layer_0[2357]; 
    assign out[5603] = layer_0[4428] & layer_0[9496]; 
    assign out[5604] = ~(layer_0[6482] | layer_0[9681]); 
    assign out[5605] = layer_0[4755] & ~layer_0[3494]; 
    assign out[5606] = layer_0[3085]; 
    assign out[5607] = ~layer_0[5773]; 
    assign out[5608] = layer_0[9883] ^ layer_0[10655]; 
    assign out[5609] = ~(layer_0[2032] | layer_0[7352]); 
    assign out[5610] = ~(layer_0[8538] ^ layer_0[2891]); 
    assign out[5611] = layer_0[6041]; 
    assign out[5612] = ~layer_0[6992]; 
    assign out[5613] = layer_0[7413]; 
    assign out[5614] = layer_0[9393] ^ layer_0[8195]; 
    assign out[5615] = layer_0[4301]; 
    assign out[5616] = layer_0[2234] ^ layer_0[8120]; 
    assign out[5617] = ~layer_0[5904]; 
    assign out[5618] = layer_0[3274]; 
    assign out[5619] = ~(layer_0[397] ^ layer_0[5587]); 
    assign out[5620] = ~(layer_0[5815] ^ layer_0[9231]); 
    assign out[5621] = ~(layer_0[7267] | layer_0[5111]); 
    assign out[5622] = layer_0[2005] & layer_0[4773]; 
    assign out[5623] = ~layer_0[2175] | (layer_0[2175] & layer_0[10785]); 
    assign out[5624] = layer_0[4535] ^ layer_0[9888]; 
    assign out[5625] = ~(layer_0[6958] ^ layer_0[8318]); 
    assign out[5626] = layer_0[6273] & ~layer_0[5191]; 
    assign out[5627] = ~layer_0[8738]; 
    assign out[5628] = ~(layer_0[54] | layer_0[4510]); 
    assign out[5629] = layer_0[4574] & layer_0[3726]; 
    assign out[5630] = ~(layer_0[10711] ^ layer_0[3488]); 
    assign out[5631] = layer_0[2509] & ~layer_0[7276]; 
    assign out[5632] = ~(layer_0[6553] | layer_0[2084]); 
    assign out[5633] = ~(layer_0[10371] ^ layer_0[460]); 
    assign out[5634] = ~layer_0[6639]; 
    assign out[5635] = layer_0[3803]; 
    assign out[5636] = layer_0[4441] & ~layer_0[615]; 
    assign out[5637] = ~(layer_0[11267] ^ layer_0[3463]); 
    assign out[5638] = layer_0[11810]; 
    assign out[5639] = ~layer_0[10281]; 
    assign out[5640] = ~(layer_0[4815] | layer_0[9698]); 
    assign out[5641] = layer_0[5151] & layer_0[9959]; 
    assign out[5642] = ~(layer_0[1687] | layer_0[2262]); 
    assign out[5643] = ~(layer_0[2163] | layer_0[8948]); 
    assign out[5644] = layer_0[10012] ^ layer_0[3945]; 
    assign out[5645] = layer_0[8682] ^ layer_0[11241]; 
    assign out[5646] = layer_0[11970]; 
    assign out[5647] = layer_0[7583]; 
    assign out[5648] = ~(layer_0[8086] ^ layer_0[10559]); 
    assign out[5649] = layer_0[8928] ^ layer_0[837]; 
    assign out[5650] = ~(layer_0[6318] ^ layer_0[382]); 
    assign out[5651] = layer_0[2531] & ~layer_0[1731]; 
    assign out[5652] = ~(layer_0[6264] ^ layer_0[10508]); 
    assign out[5653] = ~layer_0[9133] | (layer_0[9133] & layer_0[2300]); 
    assign out[5654] = layer_0[10831] & layer_0[10646]; 
    assign out[5655] = ~(layer_0[1738] | layer_0[7843]); 
    assign out[5656] = layer_0[5275] & ~layer_0[5216]; 
    assign out[5657] = layer_0[7300] ^ layer_0[10838]; 
    assign out[5658] = ~(layer_0[8699] ^ layer_0[4982]); 
    assign out[5659] = layer_0[10762] ^ layer_0[2380]; 
    assign out[5660] = layer_0[3385] & ~layer_0[10254]; 
    assign out[5661] = layer_0[3760] ^ layer_0[4076]; 
    assign out[5662] = layer_0[1899] & ~layer_0[2967]; 
    assign out[5663] = ~(layer_0[3184] ^ layer_0[311]); 
    assign out[5664] = ~layer_0[4613]; 
    assign out[5665] = ~(layer_0[4007] ^ layer_0[11580]); 
    assign out[5666] = ~(layer_0[6299] ^ layer_0[6311]); 
    assign out[5667] = layer_0[2645] ^ layer_0[6162]; 
    assign out[5668] = layer_0[241] & ~layer_0[4114]; 
    assign out[5669] = ~(layer_0[8819] | layer_0[3675]); 
    assign out[5670] = ~(layer_0[1355] | layer_0[1343]); 
    assign out[5671] = ~(layer_0[2465] | layer_0[5009]); 
    assign out[5672] = layer_0[10500] ^ layer_0[5379]; 
    assign out[5673] = ~(layer_0[7682] ^ layer_0[5428]); 
    assign out[5674] = ~layer_0[1890] | (layer_0[6389] & layer_0[1890]); 
    assign out[5675] = ~layer_0[8585] | (layer_0[8585] & layer_0[1214]); 
    assign out[5676] = layer_0[4520] & ~layer_0[7568]; 
    assign out[5677] = layer_0[5734] ^ layer_0[11646]; 
    assign out[5678] = ~layer_0[1215] | (layer_0[1215] & layer_0[1846]); 
    assign out[5679] = ~(layer_0[11231] ^ layer_0[399]); 
    assign out[5680] = layer_0[10441]; 
    assign out[5681] = layer_0[539] ^ layer_0[46]; 
    assign out[5682] = ~(layer_0[7295] | layer_0[1686]); 
    assign out[5683] = 1'b0; 
    assign out[5684] = layer_0[11437] ^ layer_0[120]; 
    assign out[5685] = layer_0[11107] ^ layer_0[1842]; 
    assign out[5686] = layer_0[9282] ^ layer_0[9555]; 
    assign out[5687] = layer_0[1288] & ~layer_0[2244]; 
    assign out[5688] = layer_0[11747] ^ layer_0[6136]; 
    assign out[5689] = ~layer_0[1270]; 
    assign out[5690] = ~layer_0[2811]; 
    assign out[5691] = ~(layer_0[6134] ^ layer_0[39]); 
    assign out[5692] = ~layer_0[1780]; 
    assign out[5693] = layer_0[10291] ^ layer_0[7051]; 
    assign out[5694] = ~(layer_0[4295] | layer_0[7360]); 
    assign out[5695] = layer_0[8004] & ~layer_0[6696]; 
    assign out[5696] = layer_0[8234] & ~layer_0[4929]; 
    assign out[5697] = layer_0[9879] ^ layer_0[828]; 
    assign out[5698] = layer_0[10037] ^ layer_0[4259]; 
    assign out[5699] = ~(layer_0[2418] ^ layer_0[1909]); 
    assign out[5700] = layer_0[6689] ^ layer_0[9648]; 
    assign out[5701] = layer_0[4098] & ~layer_0[10608]; 
    assign out[5702] = layer_0[2299] ^ layer_0[6107]; 
    assign out[5703] = ~(layer_0[7920] & layer_0[10166]); 
    assign out[5704] = ~(layer_0[4250] ^ layer_0[3312]); 
    assign out[5705] = layer_0[9135] & layer_0[7432]; 
    assign out[5706] = ~(layer_0[9001] | layer_0[5614]); 
    assign out[5707] = layer_0[5559] & ~layer_0[11120]; 
    assign out[5708] = ~layer_0[315]; 
    assign out[5709] = ~layer_0[10478]; 
    assign out[5710] = layer_0[4548] ^ layer_0[9335]; 
    assign out[5711] = ~(layer_0[10361] ^ layer_0[3620]); 
    assign out[5712] = ~(layer_0[10298] ^ layer_0[10621]); 
    assign out[5713] = ~(layer_0[9297] & layer_0[2856]); 
    assign out[5714] = layer_0[1547] ^ layer_0[4281]; 
    assign out[5715] = layer_0[4331]; 
    assign out[5716] = layer_0[10574] ^ layer_0[11522]; 
    assign out[5717] = ~(layer_0[10713] ^ layer_0[7452]); 
    assign out[5718] = ~(layer_0[834] ^ layer_0[6028]); 
    assign out[5719] = ~(layer_0[4738] ^ layer_0[6316]); 
    assign out[5720] = ~layer_0[5986] | (layer_0[5986] & layer_0[110]); 
    assign out[5721] = layer_0[7793] ^ layer_0[11463]; 
    assign out[5722] = layer_0[11129] ^ layer_0[117]; 
    assign out[5723] = layer_0[4397]; 
    assign out[5724] = layer_0[6688] ^ layer_0[9447]; 
    assign out[5725] = ~layer_0[8307]; 
    assign out[5726] = layer_0[10881] ^ layer_0[8559]; 
    assign out[5727] = ~layer_0[8734]; 
    assign out[5728] = ~(layer_0[8498] & layer_0[2707]); 
    assign out[5729] = layer_0[7029] ^ layer_0[10300]; 
    assign out[5730] = layer_0[4897] ^ layer_0[10112]; 
    assign out[5731] = layer_0[7364] ^ layer_0[5818]; 
    assign out[5732] = ~(layer_0[7184] | layer_0[7992]); 
    assign out[5733] = ~(layer_0[2527] ^ layer_0[4145]); 
    assign out[5734] = ~layer_0[8847] | (layer_0[9715] & layer_0[8847]); 
    assign out[5735] = layer_0[1044] & ~layer_0[5888]; 
    assign out[5736] = ~layer_0[871]; 
    assign out[5737] = layer_0[4455] ^ layer_0[5044]; 
    assign out[5738] = ~(layer_0[11462] | layer_0[5033]); 
    assign out[5739] = layer_0[9191] ^ layer_0[6763]; 
    assign out[5740] = ~layer_0[4997]; 
    assign out[5741] = ~layer_0[9560] | (layer_0[4041] & layer_0[9560]); 
    assign out[5742] = ~layer_0[10431]; 
    assign out[5743] = layer_0[143] ^ layer_0[8201]; 
    assign out[5744] = layer_0[681] ^ layer_0[8283]; 
    assign out[5745] = ~(layer_0[2370] | layer_0[3577]); 
    assign out[5746] = ~layer_0[11012]; 
    assign out[5747] = layer_0[6728] & ~layer_0[4234]; 
    assign out[5748] = ~layer_0[4272]; 
    assign out[5749] = layer_0[6846] & ~layer_0[2279]; 
    assign out[5750] = layer_0[8216] | layer_0[8199]; 
    assign out[5751] = layer_0[10501]; 
    assign out[5752] = ~layer_0[99]; 
    assign out[5753] = layer_0[6921] & layer_0[793]; 
    assign out[5754] = ~layer_0[7925]; 
    assign out[5755] = layer_0[8031] ^ layer_0[2468]; 
    assign out[5756] = ~(layer_0[3457] | layer_0[7703]); 
    assign out[5757] = layer_0[6540] & ~layer_0[6075]; 
    assign out[5758] = layer_0[10934]; 
    assign out[5759] = layer_0[1995] & ~layer_0[2436]; 
    assign out[5760] = ~layer_0[10961] | (layer_0[11420] & layer_0[10961]); 
    assign out[5761] = layer_0[7400] ^ layer_0[839]; 
    assign out[5762] = ~(layer_0[7979] | layer_0[730]); 
    assign out[5763] = ~layer_0[3794]; 
    assign out[5764] = layer_0[5991] ^ layer_0[11943]; 
    assign out[5765] = layer_0[6772] | layer_0[10035]; 
    assign out[5766] = layer_0[2205] ^ layer_0[3943]; 
    assign out[5767] = layer_0[3110] & ~layer_0[6411]; 
    assign out[5768] = layer_0[5853] & layer_0[9491]; 
    assign out[5769] = layer_0[3114] ^ layer_0[6632]; 
    assign out[5770] = ~(layer_0[10977] ^ layer_0[8022]); 
    assign out[5771] = layer_0[9669] ^ layer_0[3675]; 
    assign out[5772] = layer_0[290]; 
    assign out[5773] = ~(layer_0[2665] ^ layer_0[9453]); 
    assign out[5774] = layer_0[3556] ^ layer_0[5280]; 
    assign out[5775] = layer_0[5879] & ~layer_0[907]; 
    assign out[5776] = layer_0[1653] ^ layer_0[4828]; 
    assign out[5777] = ~(layer_0[5450] ^ layer_0[11630]); 
    assign out[5778] = ~layer_0[5628] | (layer_0[9730] & layer_0[5628]); 
    assign out[5779] = layer_0[8638] ^ layer_0[5451]; 
    assign out[5780] = layer_0[6872] ^ layer_0[10214]; 
    assign out[5781] = layer_0[9649] & ~layer_0[7453]; 
    assign out[5782] = layer_0[9368] & ~layer_0[8820]; 
    assign out[5783] = ~(layer_0[1310] ^ layer_0[583]); 
    assign out[5784] = layer_0[3429] & ~layer_0[11486]; 
    assign out[5785] = ~(layer_0[4953] ^ layer_0[282]); 
    assign out[5786] = layer_0[10139] ^ layer_0[1213]; 
    assign out[5787] = layer_0[9083] & ~layer_0[10159]; 
    assign out[5788] = ~layer_0[5713]; 
    assign out[5789] = layer_0[482]; 
    assign out[5790] = layer_0[11643] ^ layer_0[2725]; 
    assign out[5791] = ~(layer_0[763] ^ layer_0[1851]); 
    assign out[5792] = ~layer_0[2690]; 
    assign out[5793] = ~layer_0[425]; 
    assign out[5794] = layer_0[9498] ^ layer_0[1667]; 
    assign out[5795] = 1'b0; 
    assign out[5796] = layer_0[11326] & ~layer_0[6489]; 
    assign out[5797] = layer_0[7670] ^ layer_0[3776]; 
    assign out[5798] = ~(layer_0[4312] ^ layer_0[1350]); 
    assign out[5799] = layer_0[9215] & ~layer_0[11335]; 
    assign out[5800] = layer_0[2199] | layer_0[4208]; 
    assign out[5801] = layer_0[3126] ^ layer_0[8453]; 
    assign out[5802] = layer_0[10449] & ~layer_0[4614]; 
    assign out[5803] = layer_0[2454] & layer_0[8111]; 
    assign out[5804] = layer_0[342]; 
    assign out[5805] = ~(layer_0[7219] ^ layer_0[7405]); 
    assign out[5806] = layer_0[6884] & ~layer_0[3863]; 
    assign out[5807] = layer_0[470] ^ layer_0[4626]; 
    assign out[5808] = ~(layer_0[128] | layer_0[9668]); 
    assign out[5809] = layer_0[4909] ^ layer_0[5980]; 
    assign out[5810] = ~(layer_0[11557] | layer_0[6195]); 
    assign out[5811] = layer_0[926] & layer_0[11818]; 
    assign out[5812] = layer_0[3578] & layer_0[6476]; 
    assign out[5813] = layer_0[11431] & ~layer_0[2134]; 
    assign out[5814] = layer_0[3120] & ~layer_0[7135]; 
    assign out[5815] = layer_0[483] & ~layer_0[6175]; 
    assign out[5816] = layer_0[1495] & ~layer_0[4427]; 
    assign out[5817] = layer_0[3230] | layer_0[3127]; 
    assign out[5818] = layer_0[1568]; 
    assign out[5819] = layer_0[9793] & ~layer_0[3153]; 
    assign out[5820] = ~(layer_0[4157] & layer_0[9131]); 
    assign out[5821] = layer_0[8490] ^ layer_0[9978]; 
    assign out[5822] = ~(layer_0[9986] ^ layer_0[10296]); 
    assign out[5823] = layer_0[5382]; 
    assign out[5824] = ~layer_0[1077]; 
    assign out[5825] = layer_0[1879] ^ layer_0[5174]; 
    assign out[5826] = layer_0[7635] ^ layer_0[3128]; 
    assign out[5827] = layer_0[1412] & ~layer_0[11068]; 
    assign out[5828] = layer_0[289] ^ layer_0[4383]; 
    assign out[5829] = ~layer_0[226]; 
    assign out[5830] = layer_0[8978] & ~layer_0[3922]; 
    assign out[5831] = ~layer_0[2841]; 
    assign out[5832] = ~layer_0[3308]; 
    assign out[5833] = ~(layer_0[3311] ^ layer_0[7011]); 
    assign out[5834] = ~(layer_0[9060] ^ layer_0[7408]); 
    assign out[5835] = ~(layer_0[9214] ^ layer_0[6926]); 
    assign out[5836] = layer_0[11718] ^ layer_0[6013]; 
    assign out[5837] = ~(layer_0[3749] | layer_0[3262]); 
    assign out[5838] = ~(layer_0[8399] | layer_0[4411]); 
    assign out[5839] = layer_0[8721] ^ layer_0[2830]; 
    assign out[5840] = layer_0[4889] ^ layer_0[10335]; 
    assign out[5841] = layer_0[724] ^ layer_0[9985]; 
    assign out[5842] = layer_0[986] | layer_0[8146]; 
    assign out[5843] = layer_0[3452] ^ layer_0[7742]; 
    assign out[5844] = layer_0[7908]; 
    assign out[5845] = layer_0[694] ^ layer_0[1600]; 
    assign out[5846] = layer_0[1810] ^ layer_0[6519]; 
    assign out[5847] = layer_0[5669] & ~layer_0[4726]; 
    assign out[5848] = ~layer_0[4586] | (layer_0[9501] & layer_0[4586]); 
    assign out[5849] = layer_0[3228]; 
    assign out[5850] = layer_0[2959] & ~layer_0[2334]; 
    assign out[5851] = ~(layer_0[6906] ^ layer_0[4610]); 
    assign out[5852] = layer_0[481] & layer_0[5977]; 
    assign out[5853] = layer_0[6391] & ~layer_0[97]; 
    assign out[5854] = layer_0[237] & ~layer_0[4568]; 
    assign out[5855] = layer_0[10386] & layer_0[3694]; 
    assign out[5856] = ~(layer_0[7894] ^ layer_0[11789]); 
    assign out[5857] = layer_0[3005] & ~layer_0[6864]; 
    assign out[5858] = layer_0[6610]; 
    assign out[5859] = layer_0[8569] & ~layer_0[9745]; 
    assign out[5860] = layer_0[247] & layer_0[6783]; 
    assign out[5861] = layer_0[5102] ^ layer_0[7707]; 
    assign out[5862] = layer_0[10398] ^ layer_0[6332]; 
    assign out[5863] = ~layer_0[10177] | (layer_0[10177] & layer_0[1781]); 
    assign out[5864] = layer_0[5996] & ~layer_0[617]; 
    assign out[5865] = ~(layer_0[11475] ^ layer_0[145]); 
    assign out[5866] = ~(layer_0[2865] ^ layer_0[4051]); 
    assign out[5867] = ~(layer_0[1665] ^ layer_0[5864]); 
    assign out[5868] = ~(layer_0[2580] ^ layer_0[8503]); 
    assign out[5869] = layer_0[11075] & ~layer_0[3854]; 
    assign out[5870] = layer_0[262]; 
    assign out[5871] = ~(layer_0[10481] ^ layer_0[982]); 
    assign out[5872] = layer_0[9439] & layer_0[5881]; 
    assign out[5873] = ~layer_0[10277]; 
    assign out[5874] = layer_0[6910] & ~layer_0[8553]; 
    assign out[5875] = ~(layer_0[2216] ^ layer_0[2237]); 
    assign out[5876] = ~(layer_0[2241] ^ layer_0[4685]); 
    assign out[5877] = layer_0[1208] & ~layer_0[6255]; 
    assign out[5878] = layer_0[9120]; 
    assign out[5879] = ~layer_0[10953] | (layer_0[10953] & layer_0[489]); 
    assign out[5880] = layer_0[11760]; 
    assign out[5881] = ~(layer_0[2112] ^ layer_0[5966]); 
    assign out[5882] = ~layer_0[1812]; 
    assign out[5883] = layer_0[4224] & ~layer_0[11965]; 
    assign out[5884] = ~layer_0[6668]; 
    assign out[5885] = ~(layer_0[93] | layer_0[8160]); 
    assign out[5886] = layer_0[10185] ^ layer_0[10722]; 
    assign out[5887] = ~(layer_0[3083] ^ layer_0[964]); 
    assign out[5888] = layer_0[9228] & ~layer_0[11805]; 
    assign out[5889] = layer_0[7342] ^ layer_0[971]; 
    assign out[5890] = ~(layer_0[3191] | layer_0[1473]); 
    assign out[5891] = layer_0[2202] | layer_0[9168]; 
    assign out[5892] = layer_0[7826] & ~layer_0[3109]; 
    assign out[5893] = ~(layer_0[11681] ^ layer_0[10084]); 
    assign out[5894] = layer_0[10814]; 
    assign out[5895] = layer_0[2452] ^ layer_0[10821]; 
    assign out[5896] = ~(layer_0[2495] | layer_0[3477]); 
    assign out[5897] = ~layer_0[7804]; 
    assign out[5898] = ~(layer_0[1913] | layer_0[832]); 
    assign out[5899] = layer_0[8716]; 
    assign out[5900] = ~(layer_0[11120] ^ layer_0[4062]); 
    assign out[5901] = ~(layer_0[8739] | layer_0[4772]); 
    assign out[5902] = ~(layer_0[28] ^ layer_0[10858]); 
    assign out[5903] = layer_0[1644] & ~layer_0[3553]; 
    assign out[5904] = layer_0[7264] & ~layer_0[4308]; 
    assign out[5905] = layer_0[4557] | layer_0[10237]; 
    assign out[5906] = ~layer_0[9003]; 
    assign out[5907] = layer_0[1924]; 
    assign out[5908] = ~(layer_0[2346] & layer_0[783]); 
    assign out[5909] = ~(layer_0[2863] ^ layer_0[6150]); 
    assign out[5910] = layer_0[1800] ^ layer_0[2455]; 
    assign out[5911] = ~layer_0[9309] | (layer_0[3662] & layer_0[9309]); 
    assign out[5912] = layer_0[3204] ^ layer_0[9649]; 
    assign out[5913] = layer_0[7170] & ~layer_0[1203]; 
    assign out[5914] = layer_0[6241] | layer_0[9895]; 
    assign out[5915] = ~(layer_0[10597] | layer_0[9263]); 
    assign out[5916] = layer_0[4353] | layer_0[3481]; 
    assign out[5917] = ~layer_0[5495]; 
    assign out[5918] = ~layer_0[11421]; 
    assign out[5919] = ~(layer_0[10320] ^ layer_0[10434]); 
    assign out[5920] = layer_0[9525] & layer_0[7986]; 
    assign out[5921] = ~(layer_0[6808] | layer_0[6208]); 
    assign out[5922] = layer_0[9287] | layer_0[2459]; 
    assign out[5923] = ~layer_0[1968] | (layer_0[1968] & layer_0[2255]); 
    assign out[5924] = layer_0[5819] & ~layer_0[9507]; 
    assign out[5925] = layer_0[2708] & ~layer_0[632]; 
    assign out[5926] = layer_0[11192] & ~layer_0[1326]; 
    assign out[5927] = layer_0[11524]; 
    assign out[5928] = layer_0[5108] & ~layer_0[8697]; 
    assign out[5929] = ~layer_0[10301] | (layer_0[10301] & layer_0[5089]); 
    assign out[5930] = ~(layer_0[6808] ^ layer_0[7165]); 
    assign out[5931] = ~(layer_0[10596] ^ layer_0[8116]); 
    assign out[5932] = layer_0[9100] & layer_0[5281]; 
    assign out[5933] = ~(layer_0[6005] | layer_0[3406]); 
    assign out[5934] = layer_0[8100] ^ layer_0[3874]; 
    assign out[5935] = ~(layer_0[4778] ^ layer_0[7119]); 
    assign out[5936] = layer_0[7072] & ~layer_0[2385]; 
    assign out[5937] = ~layer_0[4973]; 
    assign out[5938] = ~(layer_0[4506] ^ layer_0[10476]); 
    assign out[5939] = ~(layer_0[7522] ^ layer_0[8938]); 
    assign out[5940] = layer_0[11316] ^ layer_0[11828]; 
    assign out[5941] = layer_0[9385]; 
    assign out[5942] = layer_0[6565] & ~layer_0[2384]; 
    assign out[5943] = ~(layer_0[11270] | layer_0[6533]); 
    assign out[5944] = layer_0[11731] ^ layer_0[3947]; 
    assign out[5945] = layer_0[4206] ^ layer_0[3967]; 
    assign out[5946] = layer_0[8830] & ~layer_0[3241]; 
    assign out[5947] = layer_0[9213]; 
    assign out[5948] = layer_0[1953] ^ layer_0[3785]; 
    assign out[5949] = layer_0[10459]; 
    assign out[5950] = ~layer_0[617]; 
    assign out[5951] = layer_0[8264] & ~layer_0[1708]; 
    assign out[5952] = ~layer_0[5958] | (layer_0[7102] & layer_0[5958]); 
    assign out[5953] = layer_0[6641] ^ layer_0[5963]; 
    assign out[5954] = layer_0[10456]; 
    assign out[5955] = layer_0[2251] ^ layer_0[1917]; 
    assign out[5956] = layer_0[530] & ~layer_0[452]; 
    assign out[5957] = layer_0[2337] ^ layer_0[10395]; 
    assign out[5958] = layer_0[5673] & ~layer_0[4956]; 
    assign out[5959] = ~(layer_0[2743] ^ layer_0[7720]); 
    assign out[5960] = layer_0[5434] ^ layer_0[1160]; 
    assign out[5961] = ~(layer_0[1190] ^ layer_0[4720]); 
    assign out[5962] = layer_0[7454] & ~layer_0[6403]; 
    assign out[5963] = layer_0[10757] & ~layer_0[7083]; 
    assign out[5964] = layer_0[5066] ^ layer_0[5070]; 
    assign out[5965] = ~layer_0[11149]; 
    assign out[5966] = ~(layer_0[1706] | layer_0[1140]); 
    assign out[5967] = layer_0[3491] & ~layer_0[9570]; 
    assign out[5968] = ~layer_0[10243]; 
    assign out[5969] = layer_0[643] & ~layer_0[7703]; 
    assign out[5970] = layer_0[420] ^ layer_0[1489]; 
    assign out[5971] = ~layer_0[5713]; 
    assign out[5972] = layer_0[8642] ^ layer_0[3797]; 
    assign out[5973] = layer_0[7226] ^ layer_0[2159]; 
    assign out[5974] = layer_0[4954] & ~layer_0[11396]; 
    assign out[5975] = layer_0[2272] ^ layer_0[10921]; 
    assign out[5976] = layer_0[6114] & ~layer_0[11661]; 
    assign out[5977] = layer_0[2191]; 
    assign out[5978] = layer_0[9958]; 
    assign out[5979] = ~layer_0[9529] | (layer_0[2458] & layer_0[9529]); 
    assign out[5980] = layer_0[3647]; 
    assign out[5981] = layer_0[11856] & ~layer_0[10397]; 
    assign out[5982] = layer_0[4097] ^ layer_0[3068]; 
    assign out[5983] = layer_0[4605] | layer_0[11464]; 
    assign out[5984] = layer_0[1664]; 
    assign out[5985] = ~(layer_0[10385] ^ layer_0[11831]); 
    assign out[5986] = ~(layer_0[467] ^ layer_0[5408]); 
    assign out[5987] = ~(layer_0[7547] ^ layer_0[527]); 
    assign out[5988] = layer_0[8670]; 
    assign out[5989] = ~(layer_0[4608] ^ layer_0[142]); 
    assign out[5990] = layer_0[8603] & layer_0[6309]; 
    assign out[5991] = layer_0[7338] ^ layer_0[3890]; 
    assign out[5992] = ~layer_0[1041]; 
    assign out[5993] = ~(layer_0[10505] ^ layer_0[849]); 
    assign out[5994] = ~(layer_0[10281] | layer_0[6365]); 
    assign out[5995] = ~(layer_0[7909] ^ layer_0[2296]); 
    assign out[5996] = layer_0[5774] ^ layer_0[1436]; 
    assign out[5997] = ~(layer_0[11238] ^ layer_0[7836]); 
    assign out[5998] = layer_0[6735] ^ layer_0[5322]; 
    assign out[5999] = ~(layer_0[8857] ^ layer_0[8994]); 
    assign out[6000] = layer_0[6812] ^ layer_0[4456]; 
    assign out[6001] = layer_0[5360]; 
    assign out[6002] = layer_0[1270] ^ layer_0[7999]; 
    assign out[6003] = layer_0[11559] ^ layer_0[1185]; 
    assign out[6004] = ~(layer_0[1773] ^ layer_0[10170]); 
    assign out[6005] = layer_0[11075] ^ layer_0[9254]; 
    assign out[6006] = layer_0[10980] & ~layer_0[10911]; 
    assign out[6007] = layer_0[7509] ^ layer_0[10493]; 
    assign out[6008] = layer_0[5966] ^ layer_0[7015]; 
    assign out[6009] = layer_0[3717] & layer_0[11473]; 
    assign out[6010] = layer_0[3373] & ~layer_0[5475]; 
    assign out[6011] = layer_0[9] ^ layer_0[9805]; 
    assign out[6012] = ~layer_0[3725]; 
    assign out[6013] = layer_0[10078] ^ layer_0[7933]; 
    assign out[6014] = ~(layer_0[5727] & layer_0[8174]); 
    assign out[6015] = layer_0[10055] ^ layer_0[4752]; 
    assign out[6016] = ~layer_0[4952]; 
    assign out[6017] = layer_0[2333]; 
    assign out[6018] = ~(layer_0[2720] ^ layer_0[931]); 
    assign out[6019] = layer_0[9200] & ~layer_0[9103]; 
    assign out[6020] = ~(layer_0[8155] ^ layer_0[1425]); 
    assign out[6021] = layer_0[11631] ^ layer_0[10269]; 
    assign out[6022] = layer_0[242] ^ layer_0[10034]; 
    assign out[6023] = ~(layer_0[3037] ^ layer_0[5362]); 
    assign out[6024] = ~layer_0[7811]; 
    assign out[6025] = layer_0[6966] | layer_0[4269]; 
    assign out[6026] = layer_0[7639] & layer_0[7521]; 
    assign out[6027] = layer_0[9807] & layer_0[8873]; 
    assign out[6028] = layer_0[10118]; 
    assign out[6029] = ~(layer_0[427] ^ layer_0[9240]); 
    assign out[6030] = layer_0[11822] ^ layer_0[9116]; 
    assign out[6031] = ~(layer_0[5137] | layer_0[9538]); 
    assign out[6032] = ~(layer_0[9102] ^ layer_0[3152]); 
    assign out[6033] = ~layer_0[8048]; 
    assign out[6034] = layer_0[11739] ^ layer_0[4631]; 
    assign out[6035] = layer_0[8449] | layer_0[2069]; 
    assign out[6036] = ~layer_0[6191]; 
    assign out[6037] = layer_0[7964] & ~layer_0[8766]; 
    assign out[6038] = layer_0[6059] & ~layer_0[7244]; 
    assign out[6039] = layer_0[7291] & ~layer_0[7529]; 
    assign out[6040] = layer_0[3266] ^ layer_0[744]; 
    assign out[6041] = ~layer_0[6205]; 
    assign out[6042] = layer_0[6692] ^ layer_0[3830]; 
    assign out[6043] = layer_0[11975] | layer_0[6852]; 
    assign out[6044] = layer_0[3917] & ~layer_0[1060]; 
    assign out[6045] = layer_0[10405] ^ layer_0[4482]; 
    assign out[6046] = ~(layer_0[7103] ^ layer_0[4887]); 
    assign out[6047] = ~layer_0[9424] | (layer_0[9424] & layer_0[539]); 
    assign out[6048] = ~(layer_0[3552] & layer_0[11396]); 
    assign out[6049] = layer_0[10042] & ~layer_0[4240]; 
    assign out[6050] = layer_0[10954] & ~layer_0[11824]; 
    assign out[6051] = ~(layer_0[1971] | layer_0[4159]); 
    assign out[6052] = layer_0[7186] ^ layer_0[7739]; 
    assign out[6053] = layer_0[3047] & ~layer_0[7021]; 
    assign out[6054] = ~layer_0[7078]; 
    assign out[6055] = layer_0[4946] ^ layer_0[204]; 
    assign out[6056] = layer_0[6862] ^ layer_0[9024]; 
    assign out[6057] = ~(layer_0[5203] ^ layer_0[3235]); 
    assign out[6058] = layer_0[9600] & ~layer_0[4555]; 
    assign out[6059] = layer_0[7514] ^ layer_0[8812]; 
    assign out[6060] = layer_0[10747] & layer_0[2532]; 
    assign out[6061] = ~(layer_0[1892] ^ layer_0[1432]); 
    assign out[6062] = layer_0[4084] & layer_0[9417]; 
    assign out[6063] = ~(layer_0[11550] ^ layer_0[4161]); 
    assign out[6064] = ~(layer_0[7493] & layer_0[10633]); 
    assign out[6065] = layer_0[8131] & layer_0[6165]; 
    assign out[6066] = layer_0[6071] ^ layer_0[7087]; 
    assign out[6067] = layer_0[11259] ^ layer_0[5950]; 
    assign out[6068] = ~(layer_0[8381] ^ layer_0[6471]); 
    assign out[6069] = ~layer_0[2149]; 
    assign out[6070] = layer_0[791] & ~layer_0[11157]; 
    assign out[6071] = ~(layer_0[446] ^ layer_0[1867]); 
    assign out[6072] = ~(layer_0[4094] | layer_0[11962]); 
    assign out[6073] = layer_0[2988] ^ layer_0[8928]; 
    assign out[6074] = layer_0[258] & ~layer_0[5463]; 
    assign out[6075] = layer_0[9317] & ~layer_0[9227]; 
    assign out[6076] = ~(layer_0[11199] ^ layer_0[11311]); 
    assign out[6077] = ~(layer_0[11886] & layer_0[10889]); 
    assign out[6078] = ~(layer_0[2750] & layer_0[2871]); 
    assign out[6079] = 1'b0; 
    assign out[6080] = layer_0[11637] ^ layer_0[5017]; 
    assign out[6081] = ~(layer_0[4306] ^ layer_0[11596]); 
    assign out[6082] = ~(layer_0[3827] ^ layer_0[5248]); 
    assign out[6083] = ~(layer_0[5678] ^ layer_0[6323]); 
    assign out[6084] = layer_0[7509] ^ layer_0[8080]; 
    assign out[6085] = layer_0[735] ^ layer_0[8821]; 
    assign out[6086] = layer_0[4606] ^ layer_0[5005]; 
    assign out[6087] = layer_0[5689] ^ layer_0[4283]; 
    assign out[6088] = layer_0[6049]; 
    assign out[6089] = layer_0[11834] ^ layer_0[8675]; 
    assign out[6090] = layer_0[1702] & ~layer_0[10128]; 
    assign out[6091] = layer_0[10770] & ~layer_0[9573]; 
    assign out[6092] = layer_0[10285] & ~layer_0[1306]; 
    assign out[6093] = layer_0[5937] & ~layer_0[10259]; 
    assign out[6094] = ~layer_0[3896]; 
    assign out[6095] = layer_0[4938] & layer_0[3687]; 
    assign out[6096] = layer_0[439] & layer_0[11564]; 
    assign out[6097] = layer_0[51] & ~layer_0[5279]; 
    assign out[6098] = ~(layer_0[7994] & layer_0[11305]); 
    assign out[6099] = layer_0[1207] & layer_0[1447]; 
    assign out[6100] = ~layer_0[7874]; 
    assign out[6101] = ~(layer_0[5814] ^ layer_0[7862]); 
    assign out[6102] = ~(layer_0[1922] ^ layer_0[2874]); 
    assign out[6103] = layer_0[1889]; 
    assign out[6104] = layer_0[6895] ^ layer_0[325]; 
    assign out[6105] = layer_0[6297] ^ layer_0[6269]; 
    assign out[6106] = layer_0[2719] ^ layer_0[4433]; 
    assign out[6107] = layer_0[5472] & ~layer_0[11000]; 
    assign out[6108] = layer_0[8652] ^ layer_0[4374]; 
    assign out[6109] = ~(layer_0[3875] ^ layer_0[4795]); 
    assign out[6110] = ~(layer_0[4166] ^ layer_0[4460]); 
    assign out[6111] = layer_0[3275] ^ layer_0[3328]; 
    assign out[6112] = layer_0[3371] & ~layer_0[6838]; 
    assign out[6113] = ~layer_0[4137]; 
    assign out[6114] = ~layer_0[9170] | (layer_0[10907] & layer_0[9170]); 
    assign out[6115] = layer_0[4021] ^ layer_0[4043]; 
    assign out[6116] = layer_0[2508] & ~layer_0[8019]; 
    assign out[6117] = layer_0[4337] ^ layer_0[2847]; 
    assign out[6118] = layer_0[9090] & ~layer_0[7070]; 
    assign out[6119] = layer_0[1255] ^ layer_0[6268]; 
    assign out[6120] = layer_0[3897] ^ layer_0[8641]; 
    assign out[6121] = ~(layer_0[5494] ^ layer_0[8705]); 
    assign out[6122] = ~layer_0[9812] | (layer_0[9812] & layer_0[3722]); 
    assign out[6123] = ~(layer_0[11774] | layer_0[8054]); 
    assign out[6124] = layer_0[11765] ^ layer_0[81]; 
    assign out[6125] = layer_0[10778] & ~layer_0[5323]; 
    assign out[6126] = layer_0[9486] & layer_0[10991]; 
    assign out[6127] = ~(layer_0[7131] ^ layer_0[7195]); 
    assign out[6128] = layer_0[11686]; 
    assign out[6129] = layer_0[4313] ^ layer_0[4016]; 
    assign out[6130] = ~layer_0[7369] | (layer_0[7369] & layer_0[3642]); 
    assign out[6131] = layer_0[493]; 
    assign out[6132] = layer_0[7679] & layer_0[8428]; 
    assign out[6133] = layer_0[4598] & ~layer_0[1377]; 
    assign out[6134] = layer_0[11282]; 
    assign out[6135] = ~(layer_0[10579] ^ layer_0[2527]); 
    assign out[6136] = layer_0[1183] & layer_0[4386]; 
    assign out[6137] = layer_0[2481] & ~layer_0[8247]; 
    assign out[6138] = ~layer_0[2344]; 
    assign out[6139] = layer_0[9454] | layer_0[1959]; 
    assign out[6140] = ~(layer_0[7790] | layer_0[7284]); 
    assign out[6141] = layer_0[10793] & layer_0[3006]; 
    assign out[6142] = ~(layer_0[10554] ^ layer_0[9581]); 
    assign out[6143] = ~layer_0[7753] | (layer_0[7753] & layer_0[3189]); 
    assign out[6144] = layer_0[8582] | layer_0[811]; 
    assign out[6145] = ~(layer_0[1448] ^ layer_0[8751]); 
    assign out[6146] = layer_0[7577] ^ layer_0[1661]; 
    assign out[6147] = ~layer_0[9713]; 
    assign out[6148] = layer_0[10493] & ~layer_0[1598]; 
    assign out[6149] = layer_0[10463] ^ layer_0[4330]; 
    assign out[6150] = ~layer_0[10140]; 
    assign out[6151] = layer_0[4125] & layer_0[8914]; 
    assign out[6152] = layer_0[5769] | layer_0[4091]; 
    assign out[6153] = layer_0[9672]; 
    assign out[6154] = ~layer_0[10343]; 
    assign out[6155] = layer_0[8096] & ~layer_0[9919]; 
    assign out[6156] = layer_0[10811] & layer_0[702]; 
    assign out[6157] = layer_0[4037] | layer_0[4051]; 
    assign out[6158] = ~(layer_0[9786] ^ layer_0[6822]); 
    assign out[6159] = layer_0[1792] & ~layer_0[11571]; 
    assign out[6160] = ~(layer_0[1808] ^ layer_0[7930]); 
    assign out[6161] = layer_0[10781]; 
    assign out[6162] = layer_0[11892] & ~layer_0[10842]; 
    assign out[6163] = layer_0[11206]; 
    assign out[6164] = ~(layer_0[6740] ^ layer_0[3666]); 
    assign out[6165] = ~(layer_0[10254] | layer_0[3374]); 
    assign out[6166] = layer_0[7555] ^ layer_0[5195]; 
    assign out[6167] = layer_0[4770] | layer_0[9780]; 
    assign out[6168] = layer_0[7468]; 
    assign out[6169] = 1'b0; 
    assign out[6170] = ~(layer_0[5447] ^ layer_0[5827]); 
    assign out[6171] = ~layer_0[7884]; 
    assign out[6172] = layer_0[261]; 
    assign out[6173] = layer_0[9969] & ~layer_0[2984]; 
    assign out[6174] = ~(layer_0[1790] | layer_0[8828]); 
    assign out[6175] = ~(layer_0[11689] ^ layer_0[4413]); 
    assign out[6176] = ~(layer_0[7178] | layer_0[11213]); 
    assign out[6177] = ~layer_0[3983]; 
    assign out[6178] = ~(layer_0[5646] ^ layer_0[9473]); 
    assign out[6179] = ~layer_0[3793]; 
    assign out[6180] = layer_0[9727] ^ layer_0[9661]; 
    assign out[6181] = layer_0[1258] ^ layer_0[7256]; 
    assign out[6182] = ~(layer_0[6686] | layer_0[11445]); 
    assign out[6183] = ~layer_0[9019]; 
    assign out[6184] = layer_0[1872] & layer_0[3237]; 
    assign out[6185] = ~(layer_0[2989] ^ layer_0[4121]); 
    assign out[6186] = layer_0[5741] & ~layer_0[5135]; 
    assign out[6187] = layer_0[2945] & ~layer_0[1162]; 
    assign out[6188] = layer_0[5167]; 
    assign out[6189] = layer_0[2940] ^ layer_0[9336]; 
    assign out[6190] = ~(layer_0[14] ^ layer_0[5144]); 
    assign out[6191] = layer_0[10914] & layer_0[8158]; 
    assign out[6192] = layer_0[7653]; 
    assign out[6193] = layer_0[9051] & ~layer_0[4723]; 
    assign out[6194] = ~(layer_0[2838] ^ layer_0[9300]); 
    assign out[6195] = layer_0[11694] ^ layer_0[871]; 
    assign out[6196] = layer_0[6837] & layer_0[7570]; 
    assign out[6197] = layer_0[4915] & ~layer_0[5224]; 
    assign out[6198] = layer_0[5422] ^ layer_0[2022]; 
    assign out[6199] = ~(layer_0[10648] ^ layer_0[2946]); 
    assign out[6200] = ~layer_0[11264]; 
    assign out[6201] = layer_0[11474] & ~layer_0[7035]; 
    assign out[6202] = layer_0[11578] ^ layer_0[11931]; 
    assign out[6203] = layer_0[5299]; 
    assign out[6204] = layer_0[5897] ^ layer_0[4344]; 
    assign out[6205] = layer_0[9251] & ~layer_0[8888]; 
    assign out[6206] = ~layer_0[2754] | (layer_0[844] & layer_0[2754]); 
    assign out[6207] = ~layer_0[6901]; 
    assign out[6208] = layer_0[11605] & ~layer_0[2637]; 
    assign out[6209] = layer_0[6954]; 
    assign out[6210] = layer_0[920] | layer_0[58]; 
    assign out[6211] = layer_0[8575] & ~layer_0[10645]; 
    assign out[6212] = layer_0[5404]; 
    assign out[6213] = 1'b0; 
    assign out[6214] = layer_0[4717] & ~layer_0[1121]; 
    assign out[6215] = ~(layer_0[9076] ^ layer_0[8849]); 
    assign out[6216] = layer_0[9358] ^ layer_0[6067]; 
    assign out[6217] = ~(layer_0[1847] ^ layer_0[3057]); 
    assign out[6218] = layer_0[3555]; 
    assign out[6219] = layer_0[4418] & ~layer_0[9920]; 
    assign out[6220] = layer_0[2824] ^ layer_0[5345]; 
    assign out[6221] = ~layer_0[10031]; 
    assign out[6222] = layer_0[9741] ^ layer_0[10129]; 
    assign out[6223] = ~layer_0[5934] | (layer_0[5934] & layer_0[3615]); 
    assign out[6224] = ~(layer_0[3169] ^ layer_0[10721]); 
    assign out[6225] = ~(layer_0[11945] ^ layer_0[8238]); 
    assign out[6226] = layer_0[3662] & ~layer_0[10140]; 
    assign out[6227] = layer_0[8855] ^ layer_0[7951]; 
    assign out[6228] = layer_0[9890] ^ layer_0[11051]; 
    assign out[6229] = layer_0[10043] & layer_0[5278]; 
    assign out[6230] = layer_0[11405]; 
    assign out[6231] = layer_0[3563] & ~layer_0[4672]; 
    assign out[6232] = ~layer_0[10906]; 
    assign out[6233] = layer_0[3813] | layer_0[9943]; 
    assign out[6234] = layer_0[2920]; 
    assign out[6235] = layer_0[4168] ^ layer_0[1187]; 
    assign out[6236] = layer_0[1431]; 
    assign out[6237] = ~(layer_0[2405] | layer_0[9677]); 
    assign out[6238] = layer_0[4304] ^ layer_0[259]; 
    assign out[6239] = ~(layer_0[1758] | layer_0[8558]); 
    assign out[6240] = ~(layer_0[4902] | layer_0[9000]); 
    assign out[6241] = ~(layer_0[9623] ^ layer_0[8732]); 
    assign out[6242] = ~layer_0[5138]; 
    assign out[6243] = layer_0[11887]; 
    assign out[6244] = layer_0[6741] & layer_0[8590]; 
    assign out[6245] = ~(layer_0[978] ^ layer_0[1530]); 
    assign out[6246] = layer_0[9198] ^ layer_0[6914]; 
    assign out[6247] = ~layer_0[9294]; 
    assign out[6248] = ~layer_0[3052]; 
    assign out[6249] = ~(layer_0[5677] | layer_0[2206]); 
    assign out[6250] = ~(layer_0[3899] ^ layer_0[3625]); 
    assign out[6251] = layer_0[3640] & ~layer_0[7799]; 
    assign out[6252] = ~(layer_0[11599] | layer_0[4488]); 
    assign out[6253] = layer_0[10005] ^ layer_0[3352]; 
    assign out[6254] = ~(layer_0[2666] ^ layer_0[7890]); 
    assign out[6255] = ~(layer_0[2789] ^ layer_0[594]); 
    assign out[6256] = ~layer_0[1152]; 
    assign out[6257] = layer_0[10189] & ~layer_0[10047]; 
    assign out[6258] = layer_0[5834]; 
    assign out[6259] = ~(layer_0[11653] | layer_0[8055]); 
    assign out[6260] = layer_0[11397] & ~layer_0[5416]; 
    assign out[6261] = ~(layer_0[7969] ^ layer_0[9822]); 
    assign out[6262] = ~(layer_0[2107] ^ layer_0[80]); 
    assign out[6263] = ~(layer_0[11037] | layer_0[10284]); 
    assign out[6264] = ~(layer_0[6676] ^ layer_0[949]); 
    assign out[6265] = layer_0[10028] & ~layer_0[495]; 
    assign out[6266] = layer_0[1986] ^ layer_0[8366]; 
    assign out[6267] = ~layer_0[6724]; 
    assign out[6268] = ~layer_0[2711] | (layer_0[2946] & layer_0[2711]); 
    assign out[6269] = layer_0[1519]; 
    assign out[6270] = layer_0[10086]; 
    assign out[6271] = layer_0[7581] ^ layer_0[9327]; 
    assign out[6272] = layer_0[3583] & layer_0[7518]; 
    assign out[6273] = layer_0[6587] & layer_0[6466]; 
    assign out[6274] = layer_0[11613] & ~layer_0[10835]; 
    assign out[6275] = layer_0[6257]; 
    assign out[6276] = layer_0[7924] ^ layer_0[3033]; 
    assign out[6277] = ~layer_0[10973]; 
    assign out[6278] = ~(layer_0[9223] ^ layer_0[9510]); 
    assign out[6279] = layer_0[476] ^ layer_0[892]; 
    assign out[6280] = ~layer_0[6191]; 
    assign out[6281] = ~layer_0[11750]; 
    assign out[6282] = layer_0[9915]; 
    assign out[6283] = ~layer_0[5402]; 
    assign out[6284] = layer_0[3621]; 
    assign out[6285] = layer_0[4373] & ~layer_0[10563]; 
    assign out[6286] = ~(layer_0[3672] ^ layer_0[3716]); 
    assign out[6287] = ~(layer_0[3921] ^ layer_0[10414]); 
    assign out[6288] = layer_0[8647] & ~layer_0[3223]; 
    assign out[6289] = ~(layer_0[2965] | layer_0[7764]); 
    assign out[6290] = layer_0[3235]; 
    assign out[6291] = layer_0[6994] & ~layer_0[10923]; 
    assign out[6292] = ~layer_0[6256]; 
    assign out[6293] = layer_0[7097] & ~layer_0[7390]; 
    assign out[6294] = ~layer_0[4454]; 
    assign out[6295] = ~(layer_0[7954] ^ layer_0[6379]); 
    assign out[6296] = ~(layer_0[4896] ^ layer_0[5253]); 
    assign out[6297] = ~(layer_0[8127] ^ layer_0[8626]); 
    assign out[6298] = layer_0[74]; 
    assign out[6299] = layer_0[11110] & ~layer_0[1411]; 
    assign out[6300] = layer_0[10473] & ~layer_0[2561]; 
    assign out[6301] = layer_0[4253] ^ layer_0[326]; 
    assign out[6302] = layer_0[9372] ^ layer_0[6042]; 
    assign out[6303] = layer_0[10748]; 
    assign out[6304] = layer_0[10107] & layer_0[3049]; 
    assign out[6305] = ~layer_0[11932]; 
    assign out[6306] = ~layer_0[8018] | (layer_0[3803] & layer_0[8018]); 
    assign out[6307] = ~(layer_0[4885] ^ layer_0[10349]); 
    assign out[6308] = ~(layer_0[8285] | layer_0[9423]); 
    assign out[6309] = ~(layer_0[10482] ^ layer_0[3504]); 
    assign out[6310] = ~(layer_0[6714] ^ layer_0[11350]); 
    assign out[6311] = layer_0[8054] ^ layer_0[5124]; 
    assign out[6312] = ~(layer_0[2087] | layer_0[1176]); 
    assign out[6313] = layer_0[6773] ^ layer_0[10448]; 
    assign out[6314] = ~(layer_0[2250] | layer_0[3543]); 
    assign out[6315] = ~layer_0[8133]; 
    assign out[6316] = ~(layer_0[7498] | layer_0[9617]); 
    assign out[6317] = ~(layer_0[4684] ^ layer_0[2072]); 
    assign out[6318] = layer_0[2800]; 
    assign out[6319] = layer_0[8030] & ~layer_0[10279]; 
    assign out[6320] = ~(layer_0[5219] ^ layer_0[8964]); 
    assign out[6321] = layer_0[2571] ^ layer_0[10313]; 
    assign out[6322] = ~layer_0[3183]; 
    assign out[6323] = layer_0[7206] & ~layer_0[10289]; 
    assign out[6324] = ~(layer_0[5152] ^ layer_0[5137]); 
    assign out[6325] = layer_0[891] & ~layer_0[4033]; 
    assign out[6326] = ~layer_0[9071] | (layer_0[9071] & layer_0[10753]); 
    assign out[6327] = ~layer_0[6374]; 
    assign out[6328] = layer_0[5580] ^ layer_0[10021]; 
    assign out[6329] = layer_0[5303] ^ layer_0[481]; 
    assign out[6330] = layer_0[1149]; 
    assign out[6331] = ~layer_0[11754]; 
    assign out[6332] = layer_0[9791] ^ layer_0[4197]; 
    assign out[6333] = layer_0[546] & layer_0[10440]; 
    assign out[6334] = ~(layer_0[357] ^ layer_0[5895]); 
    assign out[6335] = layer_0[9319] & ~layer_0[3643]; 
    assign out[6336] = layer_0[8038] & layer_0[11629]; 
    assign out[6337] = layer_0[5425] ^ layer_0[3052]; 
    assign out[6338] = layer_0[2161]; 
    assign out[6339] = layer_0[10496]; 
    assign out[6340] = ~layer_0[11030] | (layer_0[11030] & layer_0[3804]); 
    assign out[6341] = layer_0[8192] ^ layer_0[8418]; 
    assign out[6342] = ~(layer_0[130] | layer_0[5103]); 
    assign out[6343] = layer_0[4493] ^ layer_0[6046]; 
    assign out[6344] = layer_0[11858] & layer_0[3572]; 
    assign out[6345] = layer_0[4406] & ~layer_0[4593]; 
    assign out[6346] = layer_0[7648]; 
    assign out[6347] = layer_0[9419] ^ layer_0[524]; 
    assign out[6348] = layer_0[7285] & layer_0[7786]; 
    assign out[6349] = layer_0[5858] ^ layer_0[4904]; 
    assign out[6350] = layer_0[4760] ^ layer_0[8033]; 
    assign out[6351] = layer_0[1318]; 
    assign out[6352] = ~layer_0[8997]; 
    assign out[6353] = layer_0[9777]; 
    assign out[6354] = layer_0[2017] ^ layer_0[10340]; 
    assign out[6355] = layer_0[8894] & ~layer_0[4333]; 
    assign out[6356] = layer_0[4991] & ~layer_0[6879]; 
    assign out[6357] = layer_0[6581] ^ layer_0[7554]; 
    assign out[6358] = layer_0[9624] & ~layer_0[10471]; 
    assign out[6359] = ~(layer_0[10648] ^ layer_0[8099]); 
    assign out[6360] = ~(layer_0[5644] ^ layer_0[2267]); 
    assign out[6361] = ~layer_0[7110]; 
    assign out[6362] = layer_0[2557] ^ layer_0[3889]; 
    assign out[6363] = ~(layer_0[5564] | layer_0[1350]); 
    assign out[6364] = ~(layer_0[4157] | layer_0[1991]); 
    assign out[6365] = layer_0[1144] ^ layer_0[1594]; 
    assign out[6366] = layer_0[7335]; 
    assign out[6367] = layer_0[5983] & layer_0[5995]; 
    assign out[6368] = layer_0[4531]; 
    assign out[6369] = layer_0[8778] ^ layer_0[7279]; 
    assign out[6370] = layer_0[1674] ^ layer_0[4887]; 
    assign out[6371] = layer_0[10072]; 
    assign out[6372] = ~(layer_0[4025] ^ layer_0[1111]); 
    assign out[6373] = ~layer_0[6768]; 
    assign out[6374] = layer_0[9347] & layer_0[5133]; 
    assign out[6375] = layer_0[10649] ^ layer_0[8934]; 
    assign out[6376] = layer_0[3387] ^ layer_0[10561]; 
    assign out[6377] = layer_0[2672]; 
    assign out[6378] = ~(layer_0[1725] ^ layer_0[4686]); 
    assign out[6379] = ~layer_0[2654] | (layer_0[2331] & layer_0[2654]); 
    assign out[6380] = layer_0[8212] ^ layer_0[1926]; 
    assign out[6381] = ~(layer_0[1162] | layer_0[4082]); 
    assign out[6382] = ~layer_0[4564]; 
    assign out[6383] = layer_0[4539] ^ layer_0[8544]; 
    assign out[6384] = ~(layer_0[9110] ^ layer_0[8557]); 
    assign out[6385] = layer_0[11435] ^ layer_0[255]; 
    assign out[6386] = layer_0[10094] & ~layer_0[4082]; 
    assign out[6387] = layer_0[11329] ^ layer_0[11183]; 
    assign out[6388] = ~(layer_0[1735] ^ layer_0[4396]); 
    assign out[6389] = ~layer_0[7151] | (layer_0[7151] & layer_0[1559]); 
    assign out[6390] = layer_0[8818] ^ layer_0[7170]; 
    assign out[6391] = ~layer_0[1719]; 
    assign out[6392] = ~(layer_0[11521] ^ layer_0[5607]); 
    assign out[6393] = layer_0[1911] ^ layer_0[11893]; 
    assign out[6394] = layer_0[4680] ^ layer_0[7089]; 
    assign out[6395] = layer_0[283] ^ layer_0[4850]; 
    assign out[6396] = layer_0[5251] & layer_0[11547]; 
    assign out[6397] = ~(layer_0[8781] ^ layer_0[2838]); 
    assign out[6398] = layer_0[6275] ^ layer_0[7602]; 
    assign out[6399] = ~(layer_0[438] ^ layer_0[3817]); 
    assign out[6400] = layer_0[5729] ^ layer_0[10548]; 
    assign out[6401] = layer_0[5018] & ~layer_0[8147]; 
    assign out[6402] = layer_0[7293] & ~layer_0[501]; 
    assign out[6403] = ~(layer_0[4484] ^ layer_0[3887]); 
    assign out[6404] = layer_0[11989]; 
    assign out[6405] = ~(layer_0[3560] & layer_0[5918]); 
    assign out[6406] = ~(layer_0[6405] | layer_0[5542]); 
    assign out[6407] = layer_0[11430]; 
    assign out[6408] = ~(layer_0[9006] ^ layer_0[6856]); 
    assign out[6409] = ~(layer_0[7503] & layer_0[2607]); 
    assign out[6410] = ~layer_0[1264]; 
    assign out[6411] = layer_0[9817]; 
    assign out[6412] = layer_0[9974]; 
    assign out[6413] = layer_0[4985] | layer_0[2156]; 
    assign out[6414] = ~(layer_0[6194] ^ layer_0[519]); 
    assign out[6415] = ~layer_0[779] | (layer_0[2273] & layer_0[779]); 
    assign out[6416] = ~(layer_0[9480] & layer_0[11530]); 
    assign out[6417] = layer_0[11379] & layer_0[6346]; 
    assign out[6418] = ~layer_0[298] | (layer_0[2643] & layer_0[298]); 
    assign out[6419] = layer_0[2843] & ~layer_0[909]; 
    assign out[6420] = ~layer_0[11556]; 
    assign out[6421] = ~(layer_0[6055] ^ layer_0[498]); 
    assign out[6422] = layer_0[9699] & ~layer_0[3199]; 
    assign out[6423] = layer_0[10909] & layer_0[2056]; 
    assign out[6424] = ~(layer_0[7590] ^ layer_0[7879]); 
    assign out[6425] = layer_0[3017] ^ layer_0[6671]; 
    assign out[6426] = ~(layer_0[4819] ^ layer_0[11917]); 
    assign out[6427] = layer_0[11452]; 
    assign out[6428] = layer_0[2655] | layer_0[2419]; 
    assign out[6429] = ~layer_0[11853] | (layer_0[5132] & layer_0[11853]); 
    assign out[6430] = ~(layer_0[422] | layer_0[5063]); 
    assign out[6431] = ~layer_0[1801]; 
    assign out[6432] = ~layer_0[888]; 
    assign out[6433] = ~(layer_0[288] ^ layer_0[9122]); 
    assign out[6434] = layer_0[11212]; 
    assign out[6435] = layer_0[1916] | layer_0[3105]; 
    assign out[6436] = ~layer_0[10985] | (layer_0[10985] & layer_0[7618]); 
    assign out[6437] = ~layer_0[8295]; 
    assign out[6438] = layer_0[2965] | layer_0[7516]; 
    assign out[6439] = layer_0[11617] ^ layer_0[1116]; 
    assign out[6440] = ~(layer_0[5226] ^ layer_0[4477]); 
    assign out[6441] = layer_0[5138] & layer_0[5963]; 
    assign out[6442] = ~layer_0[9420]; 
    assign out[6443] = ~layer_0[8504]; 
    assign out[6444] = layer_0[2195] ^ layer_0[7068]; 
    assign out[6445] = ~(layer_0[6927] ^ layer_0[5188]); 
    assign out[6446] = layer_0[101]; 
    assign out[6447] = ~layer_0[6070] | (layer_0[6070] & layer_0[666]); 
    assign out[6448] = layer_0[1876] ^ layer_0[10280]; 
    assign out[6449] = ~(layer_0[7692] ^ layer_0[2092]); 
    assign out[6450] = layer_0[8496] ^ layer_0[5736]; 
    assign out[6451] = layer_0[4530] & ~layer_0[9878]; 
    assign out[6452] = layer_0[2660]; 
    assign out[6453] = ~(layer_0[11680] & layer_0[5257]); 
    assign out[6454] = ~layer_0[3905] | (layer_0[3905] & layer_0[7911]); 
    assign out[6455] = layer_0[5027] & layer_0[5214]; 
    assign out[6456] = layer_0[1007] ^ layer_0[10659]; 
    assign out[6457] = ~layer_0[1910]; 
    assign out[6458] = layer_0[11753]; 
    assign out[6459] = ~layer_0[4381]; 
    assign out[6460] = ~(layer_0[10639] ^ layer_0[10582]); 
    assign out[6461] = ~layer_0[8072] | (layer_0[449] & layer_0[8072]); 
    assign out[6462] = layer_0[1325] & ~layer_0[8227]; 
    assign out[6463] = ~layer_0[1154] | (layer_0[1154] & layer_0[5415]); 
    assign out[6464] = layer_0[3516] & ~layer_0[7134]; 
    assign out[6465] = layer_0[3882]; 
    assign out[6466] = ~(layer_0[5247] ^ layer_0[6084]); 
    assign out[6467] = layer_0[4254]; 
    assign out[6468] = ~layer_0[2293]; 
    assign out[6469] = layer_0[1236] ^ layer_0[9684]; 
    assign out[6470] = ~(layer_0[3868] ^ layer_0[7639]); 
    assign out[6471] = ~layer_0[5803]; 
    assign out[6472] = ~(layer_0[6112] ^ layer_0[9886]); 
    assign out[6473] = layer_0[4203] ^ layer_0[559]; 
    assign out[6474] = ~(layer_0[2773] & layer_0[7447]); 
    assign out[6475] = layer_0[7158] & ~layer_0[10270]; 
    assign out[6476] = ~(layer_0[6864] ^ layer_0[8937]); 
    assign out[6477] = ~(layer_0[4402] ^ layer_0[7060]); 
    assign out[6478] = layer_0[10987]; 
    assign out[6479] = ~layer_0[9298] | (layer_0[9298] & layer_0[11107]); 
    assign out[6480] = layer_0[7975] ^ layer_0[8908]; 
    assign out[6481] = ~(layer_0[7719] ^ layer_0[4226]); 
    assign out[6482] = layer_0[9817] & ~layer_0[9685]; 
    assign out[6483] = layer_0[11542]; 
    assign out[6484] = ~(layer_0[8499] ^ layer_0[8594]); 
    assign out[6485] = layer_0[5371]; 
    assign out[6486] = layer_0[5387]; 
    assign out[6487] = ~(layer_0[10117] ^ layer_0[5841]); 
    assign out[6488] = ~layer_0[10415]; 
    assign out[6489] = ~(layer_0[6673] & layer_0[6813]); 
    assign out[6490] = layer_0[9468] ^ layer_0[1923]; 
    assign out[6491] = layer_0[5913] ^ layer_0[6881]; 
    assign out[6492] = ~layer_0[1161]; 
    assign out[6493] = layer_0[7416] ^ layer_0[7667]; 
    assign out[6494] = ~layer_0[1127]; 
    assign out[6495] = ~(layer_0[216] ^ layer_0[4638]); 
    assign out[6496] = layer_0[11914] & ~layer_0[9057]; 
    assign out[6497] = layer_0[5472] ^ layer_0[8915]; 
    assign out[6498] = ~(layer_0[6737] ^ layer_0[4231]); 
    assign out[6499] = layer_0[10518] ^ layer_0[7484]; 
    assign out[6500] = ~layer_0[9416] | (layer_0[2616] & layer_0[9416]); 
    assign out[6501] = layer_0[6151] & ~layer_0[2363]; 
    assign out[6502] = ~(layer_0[4847] ^ layer_0[9674]); 
    assign out[6503] = layer_0[10408] & ~layer_0[3001]; 
    assign out[6504] = ~(layer_0[11855] ^ layer_0[10736]); 
    assign out[6505] = ~layer_0[7945]; 
    assign out[6506] = layer_0[5546] & ~layer_0[5659]; 
    assign out[6507] = layer_0[7778] ^ layer_0[10332]; 
    assign out[6508] = layer_0[4562] & ~layer_0[779]; 
    assign out[6509] = layer_0[1366]; 
    assign out[6510] = layer_0[3796] ^ layer_0[2281]; 
    assign out[6511] = ~(layer_0[3034] ^ layer_0[2127]); 
    assign out[6512] = ~(layer_0[5289] ^ layer_0[6496]); 
    assign out[6513] = ~(layer_0[3365] ^ layer_0[11868]); 
    assign out[6514] = ~layer_0[9093] | (layer_0[9093] & layer_0[11707]); 
    assign out[6515] = layer_0[141] ^ layer_0[4314]; 
    assign out[6516] = ~layer_0[10939] | (layer_0[10939] & layer_0[7802]); 
    assign out[6517] = layer_0[4159] ^ layer_0[4699]; 
    assign out[6518] = ~(layer_0[10295] ^ layer_0[10532]); 
    assign out[6519] = ~layer_0[4153] | (layer_0[4153] & layer_0[10910]); 
    assign out[6520] = layer_0[1371]; 
    assign out[6521] = layer_0[820] ^ layer_0[948]; 
    assign out[6522] = ~layer_0[6778] | (layer_0[5330] & layer_0[6778]); 
    assign out[6523] = layer_0[9150] | layer_0[10446]; 
    assign out[6524] = ~(layer_0[10039] ^ layer_0[11834]); 
    assign out[6525] = ~layer_0[3780]; 
    assign out[6526] = layer_0[396] ^ layer_0[2550]; 
    assign out[6527] = layer_0[2683] & ~layer_0[4210]; 
    assign out[6528] = ~layer_0[8621]; 
    assign out[6529] = ~layer_0[11875]; 
    assign out[6530] = layer_0[5712] ^ layer_0[5454]; 
    assign out[6531] = ~(layer_0[6022] ^ layer_0[3263]); 
    assign out[6532] = layer_0[4619] | layer_0[8992]; 
    assign out[6533] = layer_0[11097] ^ layer_0[957]; 
    assign out[6534] = layer_0[598] | layer_0[4282]; 
    assign out[6535] = ~layer_0[10587]; 
    assign out[6536] = ~layer_0[9005] | (layer_0[7882] & layer_0[9005]); 
    assign out[6537] = layer_0[4914]; 
    assign out[6538] = ~(layer_0[11127] ^ layer_0[6594]); 
    assign out[6539] = ~(layer_0[10603] ^ layer_0[6795]); 
    assign out[6540] = layer_0[6851] ^ layer_0[7815]; 
    assign out[6541] = ~(layer_0[6342] ^ layer_0[8589]); 
    assign out[6542] = layer_0[5160]; 
    assign out[6543] = layer_0[11472] & ~layer_0[10661]; 
    assign out[6544] = ~(layer_0[9706] ^ layer_0[6891]); 
    assign out[6545] = layer_0[3754] & ~layer_0[8472]; 
    assign out[6546] = ~(layer_0[4445] ^ layer_0[520]); 
    assign out[6547] = layer_0[9951] ^ layer_0[5317]; 
    assign out[6548] = layer_0[7893] ^ layer_0[2899]; 
    assign out[6549] = layer_0[4831]; 
    assign out[6550] = ~(layer_0[2954] & layer_0[3866]); 
    assign out[6551] = ~(layer_0[6082] ^ layer_0[9557]); 
    assign out[6552] = ~(layer_0[6692] ^ layer_0[9504]); 
    assign out[6553] = ~layer_0[413] | (layer_0[413] & layer_0[9582]); 
    assign out[6554] = layer_0[3537] ^ layer_0[1905]; 
    assign out[6555] = layer_0[11848] ^ layer_0[10712]; 
    assign out[6556] = ~layer_0[5073]; 
    assign out[6557] = ~layer_0[3136]; 
    assign out[6558] = ~layer_0[8328]; 
    assign out[6559] = ~layer_0[7141] | (layer_0[3527] & layer_0[7141]); 
    assign out[6560] = layer_0[4547] & ~layer_0[4836]; 
    assign out[6561] = layer_0[8071] | layer_0[3358]; 
    assign out[6562] = layer_0[1118]; 
    assign out[6563] = ~layer_0[8853] | (layer_0[9242] & layer_0[8853]); 
    assign out[6564] = layer_0[9423] ^ layer_0[6061]; 
    assign out[6565] = ~layer_0[10601] | (layer_0[7856] & layer_0[10601]); 
    assign out[6566] = ~layer_0[8269] | (layer_0[8269] & layer_0[2456]); 
    assign out[6567] = layer_0[7811] ^ layer_0[9610]; 
    assign out[6568] = layer_0[6752]; 
    assign out[6569] = layer_0[889] ^ layer_0[6993]; 
    assign out[6570] = ~layer_0[9326]; 
    assign out[6571] = ~layer_0[1740]; 
    assign out[6572] = ~(layer_0[8711] & layer_0[10850]); 
    assign out[6573] = layer_0[597] & layer_0[9158]; 
    assign out[6574] = ~(layer_0[7767] & layer_0[9797]); 
    assign out[6575] = layer_0[457]; 
    assign out[6576] = layer_0[7611] | layer_0[3451]; 
    assign out[6577] = layer_0[10324]; 
    assign out[6578] = layer_0[10027] ^ layer_0[7131]; 
    assign out[6579] = layer_0[7140] & ~layer_0[4459]; 
    assign out[6580] = layer_0[1318] ^ layer_0[5516]; 
    assign out[6581] = layer_0[2503] ^ layer_0[2634]; 
    assign out[6582] = ~layer_0[5479] | (layer_0[5479] & layer_0[6805]); 
    assign out[6583] = layer_0[6376] ^ layer_0[1231]; 
    assign out[6584] = ~layer_0[1483]; 
    assign out[6585] = ~layer_0[1033]; 
    assign out[6586] = layer_0[4027] & ~layer_0[1280]; 
    assign out[6587] = layer_0[3299] ^ layer_0[9196]; 
    assign out[6588] = layer_0[9867] & ~layer_0[5663]; 
    assign out[6589] = layer_0[4653] ^ layer_0[9806]; 
    assign out[6590] = ~layer_0[11787] | (layer_0[11787] & layer_0[6722]); 
    assign out[6591] = layer_0[2825] ^ layer_0[3614]; 
    assign out[6592] = ~layer_0[5737] | (layer_0[8551] & layer_0[5737]); 
    assign out[6593] = layer_0[258] ^ layer_0[11271]; 
    assign out[6594] = layer_0[7258] ^ layer_0[6443]; 
    assign out[6595] = ~layer_0[3059]; 
    assign out[6596] = ~(layer_0[2507] ^ layer_0[3853]); 
    assign out[6597] = ~(layer_0[2789] ^ layer_0[682]); 
    assign out[6598] = layer_0[11212] & layer_0[10146]; 
    assign out[6599] = ~layer_0[10226] | (layer_0[1272] & layer_0[10226]); 
    assign out[6600] = layer_0[2525]; 
    assign out[6601] = ~layer_0[11240] | (layer_0[6023] & layer_0[11240]); 
    assign out[6602] = layer_0[5370] & ~layer_0[5946]; 
    assign out[6603] = layer_0[2099] ^ layer_0[4122]; 
    assign out[6604] = layer_0[1479] & ~layer_0[11720]; 
    assign out[6605] = layer_0[10212] & ~layer_0[1736]; 
    assign out[6606] = layer_0[1796] ^ layer_0[8202]; 
    assign out[6607] = ~layer_0[1925] | (layer_0[11979] & layer_0[1925]); 
    assign out[6608] = layer_0[4943]; 
    assign out[6609] = ~layer_0[863] | (layer_0[863] & layer_0[5807]); 
    assign out[6610] = ~layer_0[3222]; 
    assign out[6611] = ~(layer_0[8611] ^ layer_0[161]); 
    assign out[6612] = ~(layer_0[4969] ^ layer_0[647]); 
    assign out[6613] = layer_0[2689] ^ layer_0[71]; 
    assign out[6614] = ~layer_0[11438]; 
    assign out[6615] = ~layer_0[1546]; 
    assign out[6616] = ~(layer_0[9997] ^ layer_0[3561]); 
    assign out[6617] = ~(layer_0[6139] ^ layer_0[691]); 
    assign out[6618] = ~(layer_0[1554] ^ layer_0[2287]); 
    assign out[6619] = layer_0[6550] ^ layer_0[10216]; 
    assign out[6620] = layer_0[6564] ^ layer_0[3995]; 
    assign out[6621] = layer_0[1068]; 
    assign out[6622] = layer_0[5436] ^ layer_0[8460]; 
    assign out[6623] = layer_0[7275] ^ layer_0[3326]; 
    assign out[6624] = ~(layer_0[5243] ^ layer_0[9308]); 
    assign out[6625] = ~layer_0[11883] | (layer_0[11883] & layer_0[1868]); 
    assign out[6626] = ~(layer_0[3218] ^ layer_0[4542]); 
    assign out[6627] = ~(layer_0[169] & layer_0[11568]); 
    assign out[6628] = ~(layer_0[8659] ^ layer_0[3828]); 
    assign out[6629] = ~(layer_0[1090] ^ layer_0[1741]); 
    assign out[6630] = layer_0[10189] ^ layer_0[9579]; 
    assign out[6631] = ~(layer_0[6439] ^ layer_0[963]); 
    assign out[6632] = ~(layer_0[8083] ^ layer_0[5170]); 
    assign out[6633] = layer_0[1875] | layer_0[9957]; 
    assign out[6634] = ~layer_0[191]; 
    assign out[6635] = ~(layer_0[10773] ^ layer_0[10349]); 
    assign out[6636] = ~(layer_0[9987] ^ layer_0[10342]); 
    assign out[6637] = layer_0[4023] & ~layer_0[159]; 
    assign out[6638] = ~(layer_0[11080] ^ layer_0[7245]); 
    assign out[6639] = layer_0[4560]; 
    assign out[6640] = ~(layer_0[10601] & layer_0[221]); 
    assign out[6641] = ~layer_0[8863]; 
    assign out[6642] = layer_0[3174] & layer_0[11842]; 
    assign out[6643] = layer_0[11275]; 
    assign out[6644] = layer_0[7810] ^ layer_0[37]; 
    assign out[6645] = ~(layer_0[9781] ^ layer_0[4872]); 
    assign out[6646] = layer_0[2762] ^ layer_0[634]; 
    assign out[6647] = ~(layer_0[2367] ^ layer_0[8074]); 
    assign out[6648] = layer_0[8650] & ~layer_0[11047]; 
    assign out[6649] = layer_0[2248] ^ layer_0[231]; 
    assign out[6650] = ~layer_0[8217]; 
    assign out[6651] = layer_0[9334]; 
    assign out[6652] = ~layer_0[9250]; 
    assign out[6653] = ~(layer_0[834] ^ layer_0[7927]); 
    assign out[6654] = ~(layer_0[5889] & layer_0[7833]); 
    assign out[6655] = layer_0[10164]; 
    assign out[6656] = layer_0[3792] & layer_0[6415]; 
    assign out[6657] = ~layer_0[5539] | (layer_0[1123] & layer_0[5539]); 
    assign out[6658] = ~(layer_0[1898] ^ layer_0[6013]); 
    assign out[6659] = ~(layer_0[5690] ^ layer_0[7155]); 
    assign out[6660] = ~(layer_0[6959] ^ layer_0[1502]); 
    assign out[6661] = ~layer_0[5658] | (layer_0[10246] & layer_0[5658]); 
    assign out[6662] = layer_0[9377] & ~layer_0[10741]; 
    assign out[6663] = ~layer_0[2276] | (layer_0[2276] & layer_0[2114]); 
    assign out[6664] = layer_0[11461] ^ layer_0[3841]; 
    assign out[6665] = layer_0[2269] ^ layer_0[1852]; 
    assign out[6666] = ~layer_0[3002]; 
    assign out[6667] = ~(layer_0[973] ^ layer_0[5929]); 
    assign out[6668] = layer_0[5645]; 
    assign out[6669] = ~(layer_0[4734] ^ layer_0[8163]); 
    assign out[6670] = layer_0[6976] | layer_0[879]; 
    assign out[6671] = ~(layer_0[6518] ^ layer_0[2181]); 
    assign out[6672] = layer_0[605] ^ layer_0[8818]; 
    assign out[6673] = layer_0[4042] | layer_0[8297]; 
    assign out[6674] = ~(layer_0[9430] ^ layer_0[4348]); 
    assign out[6675] = layer_0[4617] ^ layer_0[6092]; 
    assign out[6676] = layer_0[1097]; 
    assign out[6677] = layer_0[5113]; 
    assign out[6678] = layer_0[5768] ^ layer_0[3861]; 
    assign out[6679] = layer_0[11724] & layer_0[11244]; 
    assign out[6680] = ~(layer_0[7822] ^ layer_0[9536]); 
    assign out[6681] = ~layer_0[9043] | (layer_0[9043] & layer_0[1082]); 
    assign out[6682] = ~(layer_0[7599] ^ layer_0[6678]); 
    assign out[6683] = ~(layer_0[10598] ^ layer_0[484]); 
    assign out[6684] = ~layer_0[1711] | (layer_0[2608] & layer_0[1711]); 
    assign out[6685] = ~layer_0[8631]; 
    assign out[6686] = layer_0[6080] ^ layer_0[8011]; 
    assign out[6687] = ~layer_0[9891] | (layer_0[9891] & layer_0[1588]); 
    assign out[6688] = ~layer_0[3434] | (layer_0[3434] & layer_0[11482]); 
    assign out[6689] = ~(layer_0[2815] ^ layer_0[9611]); 
    assign out[6690] = layer_0[4848]; 
    assign out[6691] = ~layer_0[8430]; 
    assign out[6692] = ~(layer_0[8978] ^ layer_0[11236]); 
    assign out[6693] = layer_0[9708] ^ layer_0[6246]; 
    assign out[6694] = layer_0[7622]; 
    assign out[6695] = layer_0[11404] | layer_0[3942]; 
    assign out[6696] = ~(layer_0[4630] ^ layer_0[499]); 
    assign out[6697] = layer_0[6497]; 
    assign out[6698] = layer_0[7105] ^ layer_0[761]; 
    assign out[6699] = ~(layer_0[680] & layer_0[11553]); 
    assign out[6700] = ~(layer_0[6702] & layer_0[1680]); 
    assign out[6701] = ~(layer_0[1762] ^ layer_0[6147]); 
    assign out[6702] = ~(layer_0[11564] & layer_0[11436]); 
    assign out[6703] = ~(layer_0[8236] ^ layer_0[2324]); 
    assign out[6704] = layer_0[3398]; 
    assign out[6705] = ~layer_0[7935]; 
    assign out[6706] = ~(layer_0[4462] ^ layer_0[8087]); 
    assign out[6707] = layer_0[5652]; 
    assign out[6708] = ~layer_0[10563]; 
    assign out[6709] = ~layer_0[8969]; 
    assign out[6710] = ~(layer_0[10337] & layer_0[2172]); 
    assign out[6711] = ~layer_0[370] | (layer_0[235] & layer_0[370]); 
    assign out[6712] = ~(layer_0[5824] | layer_0[8976]); 
    assign out[6713] = layer_0[138] & layer_0[3129]; 
    assign out[6714] = ~(layer_0[3349] ^ layer_0[9054]); 
    assign out[6715] = ~(layer_0[3870] & layer_0[3591]); 
    assign out[6716] = ~(layer_0[10423] & layer_0[7379]); 
    assign out[6717] = layer_0[4724]; 
    assign out[6718] = ~(layer_0[1670] | layer_0[2770]); 
    assign out[6719] = ~layer_0[2211]; 
    assign out[6720] = ~(layer_0[9140] ^ layer_0[3490]); 
    assign out[6721] = layer_0[8118] ^ layer_0[10849]; 
    assign out[6722] = layer_0[3036] ^ layer_0[3974]; 
    assign out[6723] = layer_0[379]; 
    assign out[6724] = layer_0[1767]; 
    assign out[6725] = layer_0[1582] ^ layer_0[10552]; 
    assign out[6726] = ~(layer_0[5360] ^ layer_0[3137]); 
    assign out[6727] = layer_0[5686] ^ layer_0[2356]; 
    assign out[6728] = layer_0[600] | layer_0[6249]; 
    assign out[6729] = layer_0[7201] & layer_0[8373]; 
    assign out[6730] = ~(layer_0[6535] ^ layer_0[8081]); 
    assign out[6731] = ~(layer_0[11827] ^ layer_0[5731]); 
    assign out[6732] = layer_0[1945]; 
    assign out[6733] = ~layer_0[662]; 
    assign out[6734] = ~layer_0[6216] | (layer_0[11610] & layer_0[6216]); 
    assign out[6735] = ~(layer_0[3652] & layer_0[10166]); 
    assign out[6736] = layer_0[8370] & layer_0[8111]; 
    assign out[6737] = layer_0[6370] & ~layer_0[3531]; 
    assign out[6738] = layer_0[10379] ^ layer_0[11359]; 
    assign out[6739] = layer_0[277] ^ layer_0[5163]; 
    assign out[6740] = ~(layer_0[9652] ^ layer_0[156]); 
    assign out[6741] = layer_0[4764]; 
    assign out[6742] = layer_0[8249] ^ layer_0[8617]; 
    assign out[6743] = layer_0[1503]; 
    assign out[6744] = layer_0[6540] ^ layer_0[745]; 
    assign out[6745] = layer_0[10258]; 
    assign out[6746] = layer_0[5436] ^ layer_0[4820]; 
    assign out[6747] = layer_0[8384]; 
    assign out[6748] = ~layer_0[5007] | (layer_0[5007] & layer_0[675]); 
    assign out[6749] = layer_0[3388] ^ layer_0[6127]; 
    assign out[6750] = layer_0[10357] ^ layer_0[3811]; 
    assign out[6751] = layer_0[5135]; 
    assign out[6752] = ~(layer_0[4130] | layer_0[11746]); 
    assign out[6753] = layer_0[4811] ^ layer_0[2034]; 
    assign out[6754] = layer_0[10943]; 
    assign out[6755] = ~(layer_0[1345] ^ layer_0[7938]); 
    assign out[6756] = layer_0[7297] ^ layer_0[3711]; 
    assign out[6757] = ~(layer_0[1814] ^ layer_0[5412]); 
    assign out[6758] = layer_0[4012] | layer_0[2554]; 
    assign out[6759] = layer_0[11365] | layer_0[1929]; 
    assign out[6760] = ~(layer_0[6334] ^ layer_0[3427]); 
    assign out[6761] = ~(layer_0[8627] | layer_0[341]); 
    assign out[6762] = ~layer_0[5072]; 
    assign out[6763] = ~(layer_0[10124] ^ layer_0[61]); 
    assign out[6764] = layer_0[9896] ^ layer_0[2893]; 
    assign out[6765] = layer_0[6745] ^ layer_0[616]; 
    assign out[6766] = layer_0[3022] ^ layer_0[10319]; 
    assign out[6767] = layer_0[5508] & ~layer_0[6156]; 
    assign out[6768] = ~(layer_0[3180] ^ layer_0[6744]); 
    assign out[6769] = layer_0[10718] & ~layer_0[6537]; 
    assign out[6770] = ~layer_0[8420] | (layer_0[3378] & layer_0[8420]); 
    assign out[6771] = layer_0[5236]; 
    assign out[6772] = ~layer_0[2270]; 
    assign out[6773] = layer_0[2118] & layer_0[11913]; 
    assign out[6774] = ~(layer_0[6936] | layer_0[2692]); 
    assign out[6775] = layer_0[8975] ^ layer_0[3601]; 
    assign out[6776] = ~layer_0[1155]; 
    assign out[6777] = layer_0[3044] & ~layer_0[923]; 
    assign out[6778] = layer_0[11382] ^ layer_0[5119]; 
    assign out[6779] = layer_0[4292] ^ layer_0[6344]; 
    assign out[6780] = ~layer_0[10799]; 
    assign out[6781] = ~layer_0[4537]; 
    assign out[6782] = ~(layer_0[6124] | layer_0[983]); 
    assign out[6783] = layer_0[5965]; 
    assign out[6784] = layer_0[6868] | layer_0[11100]; 
    assign out[6785] = ~(layer_0[9058] ^ layer_0[10546]); 
    assign out[6786] = ~(layer_0[5120] ^ layer_0[5468]); 
    assign out[6787] = ~(layer_0[5054] | layer_0[11003]); 
    assign out[6788] = layer_0[11780] ^ layer_0[4742]; 
    assign out[6789] = ~layer_0[4644] | (layer_0[4321] & layer_0[4644]); 
    assign out[6790] = ~layer_0[11729]; 
    assign out[6791] = layer_0[7414] & ~layer_0[11315]; 
    assign out[6792] = ~(layer_0[10001] ^ layer_0[10290]); 
    assign out[6793] = ~layer_0[8440] | (layer_0[8680] & layer_0[8440]); 
    assign out[6794] = ~layer_0[10343] | (layer_0[856] & layer_0[10343]); 
    assign out[6795] = ~(layer_0[11241] ^ layer_0[8367]); 
    assign out[6796] = layer_0[3566] & ~layer_0[10125]; 
    assign out[6797] = ~(layer_0[9861] ^ layer_0[8195]); 
    assign out[6798] = ~(layer_0[9097] & layer_0[10665]); 
    assign out[6799] = layer_0[9790] & ~layer_0[6033]; 
    assign out[6800] = ~(layer_0[3741] ^ layer_0[10477]); 
    assign out[6801] = layer_0[11515] ^ layer_0[519]; 
    assign out[6802] = ~layer_0[741]; 
    assign out[6803] = ~layer_0[6563] | (layer_0[3481] & layer_0[6563]); 
    assign out[6804] = layer_0[5254]; 
    assign out[6805] = layer_0[10010] ^ layer_0[3759]; 
    assign out[6806] = ~(layer_0[7955] & layer_0[3318]); 
    assign out[6807] = layer_0[8905] ^ layer_0[1220]; 
    assign out[6808] = layer_0[11049] & ~layer_0[8775]; 
    assign out[6809] = layer_0[11658] & layer_0[6481]; 
    assign out[6810] = layer_0[10000]; 
    assign out[6811] = ~layer_0[10199] | (layer_0[10199] & layer_0[9527]); 
    assign out[6812] = ~layer_0[3232] | (layer_0[3232] & layer_0[2625]); 
    assign out[6813] = layer_0[8946] ^ layer_0[3475]; 
    assign out[6814] = layer_0[9140] ^ layer_0[6604]; 
    assign out[6815] = ~(layer_0[7555] ^ layer_0[5877]); 
    assign out[6816] = layer_0[536] ^ layer_0[5738]; 
    assign out[6817] = layer_0[960] & ~layer_0[11755]; 
    assign out[6818] = layer_0[5867] ^ layer_0[11576]; 
    assign out[6819] = ~(layer_0[8136] & layer_0[7494]); 
    assign out[6820] = ~layer_0[11853]; 
    assign out[6821] = ~(layer_0[4690] ^ layer_0[2323]); 
    assign out[6822] = layer_0[8493] & ~layer_0[1168]; 
    assign out[6823] = layer_0[9277] ^ layer_0[9732]; 
    assign out[6824] = ~layer_0[5730] | (layer_0[1533] & layer_0[5730]); 
    assign out[6825] = layer_0[975]; 
    assign out[6826] = layer_0[5754] & ~layer_0[1208]; 
    assign out[6827] = ~(layer_0[2981] ^ layer_0[6037]); 
    assign out[6828] = layer_0[5605] ^ layer_0[7037]; 
    assign out[6829] = layer_0[9747] ^ layer_0[6977]; 
    assign out[6830] = ~(layer_0[3898] ^ layer_0[11205]); 
    assign out[6831] = ~(layer_0[2909] ^ layer_0[7929]); 
    assign out[6832] = layer_0[3678] ^ layer_0[11089]; 
    assign out[6833] = layer_0[2536] ^ layer_0[917]; 
    assign out[6834] = ~layer_0[3695] | (layer_0[514] & layer_0[3695]); 
    assign out[6835] = ~(layer_0[8094] ^ layer_0[7596]); 
    assign out[6836] = layer_0[5021]; 
    assign out[6837] = ~layer_0[2266]; 
    assign out[6838] = ~(layer_0[638] ^ layer_0[10847]); 
    assign out[6839] = ~(layer_0[32] & layer_0[10438]); 
    assign out[6840] = layer_0[4640] ^ layer_0[7535]; 
    assign out[6841] = layer_0[5221]; 
    assign out[6842] = ~layer_0[7156]; 
    assign out[6843] = layer_0[1772] ^ layer_0[8725]; 
    assign out[6844] = layer_0[1717] & ~layer_0[6181]; 
    assign out[6845] = ~(layer_0[882] ^ layer_0[10060]); 
    assign out[6846] = layer_0[2136] ^ layer_0[9035]; 
    assign out[6847] = ~layer_0[7770]; 
    assign out[6848] = ~(layer_0[717] ^ layer_0[7995]); 
    assign out[6849] = layer_0[7628] & layer_0[10889]; 
    assign out[6850] = layer_0[2228] ^ layer_0[1543]; 
    assign out[6851] = ~(layer_0[8636] ^ layer_0[2541]); 
    assign out[6852] = ~(layer_0[7860] ^ layer_0[5232]); 
    assign out[6853] = ~(layer_0[1022] ^ layer_0[3773]); 
    assign out[6854] = layer_0[5500]; 
    assign out[6855] = ~(layer_0[2457] & layer_0[1317]); 
    assign out[6856] = ~(layer_0[465] & layer_0[9245]); 
    assign out[6857] = ~(layer_0[6633] ^ layer_0[967]); 
    assign out[6858] = ~layer_0[8194] | (layer_0[8194] & layer_0[3337]); 
    assign out[6859] = layer_0[9353] ^ layer_0[7736]; 
    assign out[6860] = layer_0[3872] ^ layer_0[3269]; 
    assign out[6861] = layer_0[7444] ^ layer_0[10136]; 
    assign out[6862] = layer_0[4637] | layer_0[11131]; 
    assign out[6863] = ~(layer_0[302] ^ layer_0[9889]); 
    assign out[6864] = layer_0[1930] | layer_0[6293]; 
    assign out[6865] = layer_0[11997]; 
    assign out[6866] = ~(layer_0[8137] ^ layer_0[8497]); 
    assign out[6867] = ~layer_0[5052] | (layer_0[6225] & layer_0[5052]); 
    assign out[6868] = layer_0[2980] ^ layer_0[8703]; 
    assign out[6869] = ~(layer_0[4808] ^ layer_0[6375]); 
    assign out[6870] = ~(layer_0[7005] ^ layer_0[327]); 
    assign out[6871] = ~layer_0[609] | (layer_0[609] & layer_0[3251]); 
    assign out[6872] = ~layer_0[8924]; 
    assign out[6873] = ~(layer_0[4633] ^ layer_0[5955]); 
    assign out[6874] = ~layer_0[8431] | (layer_0[8339] & layer_0[8431]); 
    assign out[6875] = layer_0[7434] & layer_0[1232]; 
    assign out[6876] = layer_0[2046] & ~layer_0[4336]; 
    assign out[6877] = ~(layer_0[9294] ^ layer_0[9142]); 
    assign out[6878] = ~layer_0[5924]; 
    assign out[6879] = layer_0[4517] | layer_0[2115]; 
    assign out[6880] = layer_0[6462] ^ layer_0[10880]; 
    assign out[6881] = layer_0[9160] ^ layer_0[21]; 
    assign out[6882] = ~(layer_0[8875] & layer_0[6259]); 
    assign out[6883] = ~layer_0[8731] | (layer_0[6598] & layer_0[8731]); 
    assign out[6884] = layer_0[8907] ^ layer_0[7866]; 
    assign out[6885] = ~layer_0[8581] | (layer_0[9802] & layer_0[8581]); 
    assign out[6886] = ~layer_0[11920]; 
    assign out[6887] = layer_0[2907] ^ layer_0[8679]; 
    assign out[6888] = layer_0[7331] ^ layer_0[2467]; 
    assign out[6889] = ~(layer_0[3020] | layer_0[10852]); 
    assign out[6890] = layer_0[8637]; 
    assign out[6891] = ~(layer_0[1957] ^ layer_0[11672]); 
    assign out[6892] = ~layer_0[11957]; 
    assign out[6893] = ~(layer_0[9991] & layer_0[3371]); 
    assign out[6894] = ~(layer_0[7391] | layer_0[11344]); 
    assign out[6895] = layer_0[2572] ^ layer_0[2090]; 
    assign out[6896] = layer_0[7255] & ~layer_0[8307]; 
    assign out[6897] = layer_0[6438]; 
    assign out[6898] = ~(layer_0[2702] ^ layer_0[1323]); 
    assign out[6899] = ~layer_0[3265]; 
    assign out[6900] = ~(layer_0[9246] ^ layer_0[3635]); 
    assign out[6901] = layer_0[10005] ^ layer_0[387]; 
    assign out[6902] = layer_0[4492] | layer_0[7527]; 
    assign out[6903] = layer_0[2849] ^ layer_0[3333]; 
    assign out[6904] = layer_0[11297] ^ layer_0[2323]; 
    assign out[6905] = layer_0[10006] | layer_0[3453]; 
    assign out[6906] = ~(layer_0[10938] ^ layer_0[442]); 
    assign out[6907] = layer_0[7026] ^ layer_0[942]; 
    assign out[6908] = layer_0[11103]; 
    assign out[6909] = ~layer_0[1348] | (layer_0[10844] & layer_0[1348]); 
    assign out[6910] = ~layer_0[3660]; 
    assign out[6911] = layer_0[3291] ^ layer_0[8228]; 
    assign out[6912] = layer_0[11540] ^ layer_0[5413]; 
    assign out[6913] = layer_0[7752] & layer_0[8753]; 
    assign out[6914] = layer_0[1649] ^ layer_0[5573]; 
    assign out[6915] = layer_0[9500]; 
    assign out[6916] = layer_0[6078] | layer_0[2077]; 
    assign out[6917] = layer_0[7774] ^ layer_0[11923]; 
    assign out[6918] = ~(layer_0[3032] & layer_0[9230]); 
    assign out[6919] = layer_0[10111]; 
    assign out[6920] = layer_0[995]; 
    assign out[6921] = ~layer_0[8542]; 
    assign out[6922] = ~(layer_0[9637] ^ layer_0[6049]); 
    assign out[6923] = ~layer_0[9167]; 
    assign out[6924] = layer_0[4944]; 
    assign out[6925] = layer_0[7496] ^ layer_0[7590]; 
    assign out[6926] = ~layer_0[8328] | (layer_0[1440] & layer_0[8328]); 
    assign out[6927] = ~(layer_0[5304] & layer_0[8782]); 
    assign out[6928] = ~(layer_0[3325] ^ layer_0[4188]); 
    assign out[6929] = layer_0[8162] & layer_0[10209]; 
    assign out[6930] = layer_0[6284]; 
    assign out[6931] = ~(layer_0[5423] & layer_0[8605]); 
    assign out[6932] = layer_0[7326] & ~layer_0[10647]; 
    assign out[6933] = ~layer_0[7760]; 
    assign out[6934] = ~layer_0[9356]; 
    assign out[6935] = layer_0[184]; 
    assign out[6936] = layer_0[95] ^ layer_0[8555]; 
    assign out[6937] = ~layer_0[395]; 
    assign out[6938] = ~layer_0[8952]; 
    assign out[6939] = layer_0[1094]; 
    assign out[6940] = layer_0[6306] & ~layer_0[6967]; 
    assign out[6941] = ~layer_0[5949]; 
    assign out[6942] = layer_0[90] ^ layer_0[1975]; 
    assign out[6943] = layer_0[5410] ^ layer_0[7807]; 
    assign out[6944] = layer_0[6687]; 
    assign out[6945] = ~(layer_0[2664] ^ layer_0[7320]); 
    assign out[6946] = layer_0[4797] | layer_0[6009]; 
    assign out[6947] = layer_0[8999] ^ layer_0[11663]; 
    assign out[6948] = ~layer_0[525]; 
    assign out[6949] = ~(layer_0[1614] ^ layer_0[4303]); 
    assign out[6950] = layer_0[10331]; 
    assign out[6951] = ~(layer_0[5526] ^ layer_0[2569]); 
    assign out[6952] = ~layer_0[10125]; 
    assign out[6953] = layer_0[10119] ^ layer_0[3454]; 
    assign out[6954] = ~layer_0[8999] | (layer_0[8999] & layer_0[1153]); 
    assign out[6955] = ~(layer_0[9486] ^ layer_0[2200]); 
    assign out[6956] = layer_0[1525] ^ layer_0[9148]; 
    assign out[6957] = layer_0[4412]; 
    assign out[6958] = ~layer_0[9894] | (layer_0[1076] & layer_0[9894]); 
    assign out[6959] = ~(layer_0[11844] ^ layer_0[8270]); 
    assign out[6960] = layer_0[4278] ^ layer_0[6653]; 
    assign out[6961] = layer_0[2222] & ~layer_0[4501]; 
    assign out[6962] = layer_0[1157] ^ layer_0[6697]; 
    assign out[6963] = layer_0[6456] ^ layer_0[1802]; 
    assign out[6964] = layer_0[8784] ^ layer_0[11960]; 
    assign out[6965] = ~layer_0[6840]; 
    assign out[6966] = layer_0[9755]; 
    assign out[6967] = layer_0[2908] ^ layer_0[3605]; 
    assign out[6968] = layer_0[7096] ^ layer_0[11388]; 
    assign out[6969] = ~layer_0[5842] | (layer_0[5842] & layer_0[8314]); 
    assign out[6970] = layer_0[3904] ^ layer_0[9503]; 
    assign out[6971] = ~layer_0[3209]; 
    assign out[6972] = layer_0[181] & layer_0[6786]; 
    assign out[6973] = ~(layer_0[10606] ^ layer_0[9172]); 
    assign out[6974] = ~(layer_0[1774] ^ layer_0[7272]); 
    assign out[6975] = layer_0[8005] ^ layer_0[8424]; 
    assign out[6976] = ~layer_0[8829] | (layer_0[8829] & layer_0[4067]); 
    assign out[6977] = layer_0[3914] ^ layer_0[8206]; 
    assign out[6978] = ~(layer_0[2035] | layer_0[5848]); 
    assign out[6979] = layer_0[4373] ^ layer_0[4453]; 
    assign out[6980] = ~layer_0[8523]; 
    assign out[6981] = ~(layer_0[6493] ^ layer_0[6383]); 
    assign out[6982] = ~(layer_0[4754] ^ layer_0[1901]); 
    assign out[6983] = layer_0[2614] & ~layer_0[1965]; 
    assign out[6984] = ~(layer_0[2757] ^ layer_0[11443]); 
    assign out[6985] = ~layer_0[565] | (layer_0[5147] & layer_0[565]); 
    assign out[6986] = layer_0[10229]; 
    assign out[6987] = ~(layer_0[5700] ^ layer_0[6675]); 
    assign out[6988] = layer_0[2396] | layer_0[11639]; 
    assign out[6989] = ~(layer_0[816] ^ layer_0[10742]); 
    assign out[6990] = ~layer_0[3811] | (layer_0[3811] & layer_0[11648]); 
    assign out[6991] = ~(layer_0[8204] ^ layer_0[8224]); 
    assign out[6992] = ~(layer_0[3801] ^ layer_0[7182]); 
    assign out[6993] = layer_0[11504]; 
    assign out[6994] = layer_0[9388] ^ layer_0[829]; 
    assign out[6995] = layer_0[7311]; 
    assign out[6996] = ~layer_0[6684]; 
    assign out[6997] = layer_0[9843] ^ layer_0[4781]; 
    assign out[6998] = ~(layer_0[7070] ^ layer_0[2029]); 
    assign out[6999] = layer_0[10056] ^ layer_0[8632]; 
    assign out[7000] = layer_0[8763] & layer_0[11456]; 
    assign out[7001] = ~(layer_0[819] | layer_0[1912]); 
    assign out[7002] = ~(layer_0[3292] & layer_0[5459]); 
    assign out[7003] = layer_0[650]; 
    assign out[7004] = ~layer_0[2378]; 
    assign out[7005] = layer_0[8129] ^ layer_0[5999]; 
    assign out[7006] = layer_0[9073] & layer_0[10761]; 
    assign out[7007] = layer_0[4831] ^ layer_0[822]; 
    assign out[7008] = layer_0[2198] ^ layer_0[10017]; 
    assign out[7009] = ~(layer_0[5293] & layer_0[9963]); 
    assign out[7010] = ~layer_0[2646]; 
    assign out[7011] = layer_0[4670]; 
    assign out[7012] = layer_0[6102] ^ layer_0[10996]; 
    assign out[7013] = layer_0[11687] ^ layer_0[9041]; 
    assign out[7014] = layer_0[8242]; 
    assign out[7015] = layer_0[8838] ^ layer_0[3060]; 
    assign out[7016] = ~(layer_0[7695] ^ layer_0[3574]); 
    assign out[7017] = ~(layer_0[1177] & layer_0[8060]); 
    assign out[7018] = ~(layer_0[4003] ^ layer_0[9221]); 
    assign out[7019] = ~(layer_0[5329] ^ layer_0[5122]); 
    assign out[7020] = layer_0[3170] ^ layer_0[11348]; 
    assign out[7021] = layer_0[2633] ^ layer_0[3447]; 
    assign out[7022] = ~(layer_0[11161] ^ layer_0[9101]); 
    assign out[7023] = layer_0[5585] ^ layer_0[1018]; 
    assign out[7024] = layer_0[10762] ^ layer_0[4238]; 
    assign out[7025] = ~layer_0[182] | (layer_0[6621] & layer_0[182]); 
    assign out[7026] = ~(layer_0[5602] ^ layer_0[11531]); 
    assign out[7027] = layer_0[2031]; 
    assign out[7028] = layer_0[4100] | layer_0[7284]; 
    assign out[7029] = ~layer_0[2691]; 
    assign out[7030] = layer_0[27]; 
    assign out[7031] = layer_0[10047] & layer_0[6950]; 
    assign out[7032] = ~layer_0[2229] | (layer_0[5352] & layer_0[2229]); 
    assign out[7033] = ~(layer_0[4599] | layer_0[5300]); 
    assign out[7034] = layer_0[8303] | layer_0[1713]; 
    assign out[7035] = layer_0[412] ^ layer_0[4169]; 
    assign out[7036] = layer_0[1703] & ~layer_0[8115]; 
    assign out[7037] = layer_0[3710] ^ layer_0[9226]; 
    assign out[7038] = ~layer_0[10122]; 
    assign out[7039] = ~(layer_0[6528] | layer_0[10122]); 
    assign out[7040] = ~(layer_0[1571] | layer_0[11370]); 
    assign out[7041] = ~layer_0[8865]; 
    assign out[7042] = layer_0[1109] ^ layer_0[1799]; 
    assign out[7043] = layer_0[10300]; 
    assign out[7044] = layer_0[11945] ^ layer_0[1521]; 
    assign out[7045] = ~(layer_0[10366] & layer_0[342]); 
    assign out[7046] = layer_0[3855] ^ layer_0[6182]; 
    assign out[7047] = layer_0[8991]; 
    assign out[7048] = ~layer_0[5312]; 
    assign out[7049] = ~layer_0[883]; 
    assign out[7050] = ~(layer_0[10938] & layer_0[9716]); 
    assign out[7051] = ~(layer_0[11573] ^ layer_0[3147]); 
    assign out[7052] = ~layer_0[114] | (layer_0[8471] & layer_0[114]); 
    assign out[7053] = ~(layer_0[3176] & layer_0[7109]); 
    assign out[7054] = layer_0[11822]; 
    assign out[7055] = ~(layer_0[9273] ^ layer_0[8916]); 
    assign out[7056] = layer_0[2627] ^ layer_0[2974]; 
    assign out[7057] = layer_0[1900]; 
    assign out[7058] = ~(layer_0[2732] ^ layer_0[2296]); 
    assign out[7059] = layer_0[2221] & ~layer_0[3384]; 
    assign out[7060] = layer_0[772] ^ layer_0[1115]; 
    assign out[7061] = ~(layer_0[1745] & layer_0[9591]); 
    assign out[7062] = ~layer_0[9106]; 
    assign out[7063] = layer_0[3405] ^ layer_0[1635]; 
    assign out[7064] = layer_0[1647] ^ layer_0[132]; 
    assign out[7065] = layer_0[10744] ^ layer_0[4801]; 
    assign out[7066] = layer_0[3103]; 
    assign out[7067] = layer_0[10573] ^ layer_0[6787]; 
    assign out[7068] = layer_0[5171]; 
    assign out[7069] = ~layer_0[408] | (layer_0[7079] & layer_0[408]); 
    assign out[7070] = layer_0[11706] & layer_0[765]; 
    assign out[7071] = layer_0[5987] ^ layer_0[7844]; 
    assign out[7072] = layer_0[1744]; 
    assign out[7073] = ~layer_0[339] | (layer_0[339] & layer_0[5439]); 
    assign out[7074] = ~layer_0[3611]; 
    assign out[7075] = layer_0[8908]; 
    assign out[7076] = layer_0[3621] ^ layer_0[6086]; 
    assign out[7077] = ~(layer_0[9572] ^ layer_0[11835]); 
    assign out[7078] = layer_0[10840] ^ layer_0[7998]; 
    assign out[7079] = layer_0[1298] ^ layer_0[1664]; 
    assign out[7080] = layer_0[10690] ^ layer_0[4784]; 
    assign out[7081] = ~layer_0[7319] | (layer_0[7319] & layer_0[1245]); 
    assign out[7082] = ~(layer_0[10801] ^ layer_0[5344]); 
    assign out[7083] = layer_0[5157] & ~layer_0[1675]; 
    assign out[7084] = ~layer_0[4042] | (layer_0[4042] & layer_0[10457]); 
    assign out[7085] = layer_0[1867] ^ layer_0[5140]; 
    assign out[7086] = ~(layer_0[2698] & layer_0[11867]); 
    assign out[7087] = ~layer_0[9940]; 
    assign out[7088] = layer_0[3159] | layer_0[4785]; 
    assign out[7089] = layer_0[11922]; 
    assign out[7090] = layer_0[1012]; 
    assign out[7091] = ~layer_0[9039] | (layer_0[9039] & layer_0[954]); 
    assign out[7092] = layer_0[2624] ^ layer_0[4354]; 
    assign out[7093] = layer_0[9547] & ~layer_0[1950]; 
    assign out[7094] = ~layer_0[6730]; 
    assign out[7095] = ~(layer_0[19] ^ layer_0[508]); 
    assign out[7096] = ~(layer_0[7406] ^ layer_0[11054]); 
    assign out[7097] = ~layer_0[5120]; 
    assign out[7098] = layer_0[7899] | layer_0[139]; 
    assign out[7099] = ~layer_0[6324] | (layer_0[1272] & layer_0[6324]); 
    assign out[7100] = layer_0[9070]; 
    assign out[7101] = ~layer_0[1739] | (layer_0[1739] & layer_0[9712]); 
    assign out[7102] = layer_0[8749] ^ layer_0[2861]; 
    assign out[7103] = layer_0[9098] & ~layer_0[8546]; 
    assign out[7104] = ~layer_0[9004] | (layer_0[9149] & layer_0[9004]); 
    assign out[7105] = layer_0[5306] & ~layer_0[9918]; 
    assign out[7106] = layer_0[4479] ^ layer_0[9768]; 
    assign out[7107] = layer_0[4315] | layer_0[11918]; 
    assign out[7108] = ~layer_0[7367] | (layer_0[1392] & layer_0[7367]); 
    assign out[7109] = layer_0[7213] | layer_0[11433]; 
    assign out[7110] = ~layer_0[3944] | (layer_0[3944] & layer_0[10173]); 
    assign out[7111] = layer_0[7838] ^ layer_0[8075]; 
    assign out[7112] = layer_0[640]; 
    assign out[7113] = ~layer_0[6623] | (layer_0[6623] & layer_0[2934]); 
    assign out[7114] = ~(layer_0[812] & layer_0[7162]); 
    assign out[7115] = ~layer_0[8774]; 
    assign out[7116] = ~layer_0[9709] | (layer_0[9709] & layer_0[4078]); 
    assign out[7117] = ~(layer_0[347] ^ layer_0[6461]); 
    assign out[7118] = ~layer_0[11495] | (layer_0[11495] & layer_0[3404]); 
    assign out[7119] = ~(layer_0[26] ^ layer_0[1032]); 
    assign out[7120] = ~(layer_0[1861] ^ layer_0[9350]); 
    assign out[7121] = layer_0[8666] ^ layer_0[11549]; 
    assign out[7122] = layer_0[3641]; 
    assign out[7123] = ~(layer_0[1321] ^ layer_0[10695]); 
    assign out[7124] = layer_0[4384] | layer_0[2190]; 
    assign out[7125] = layer_0[8618]; 
    assign out[7126] = ~layer_0[42]; 
    assign out[7127] = layer_0[4370] ^ layer_0[291]; 
    assign out[7128] = ~(layer_0[9030] | layer_0[7384]); 
    assign out[7129] = ~layer_0[8291]; 
    assign out[7130] = ~(layer_0[7475] ^ layer_0[10013]); 
    assign out[7131] = layer_0[11414] ^ layer_0[2937]; 
    assign out[7132] = layer_0[2824]; 
    assign out[7133] = ~layer_0[5675] | (layer_0[134] & layer_0[5675]); 
    assign out[7134] = ~layer_0[5237] | (layer_0[5237] & layer_0[2071]); 
    assign out[7135] = ~(layer_0[2872] ^ layer_0[1684]); 
    assign out[7136] = layer_0[7700] ^ layer_0[2314]; 
    assign out[7137] = layer_0[8637] & layer_0[2024]; 
    assign out[7138] = ~(layer_0[7100] ^ layer_0[6089]); 
    assign out[7139] = ~(layer_0[10935] ^ layer_0[4445]); 
    assign out[7140] = layer_0[1935] ^ layer_0[11921]; 
    assign out[7141] = ~layer_0[11453]; 
    assign out[7142] = layer_0[11322] ^ layer_0[7744]; 
    assign out[7143] = ~(layer_0[10885] & layer_0[984]); 
    assign out[7144] = layer_0[1973]; 
    assign out[7145] = ~layer_0[62] | (layer_0[8413] & layer_0[62]); 
    assign out[7146] = layer_0[3651]; 
    assign out[7147] = ~(layer_0[8572] & layer_0[7959]); 
    assign out[7148] = layer_0[11916] ^ layer_0[7940]; 
    assign out[7149] = ~(layer_0[9770] & layer_0[7950]); 
    assign out[7150] = ~layer_0[2535] | (layer_0[8604] & layer_0[2535]); 
    assign out[7151] = ~layer_0[1324] | (layer_0[1324] & layer_0[848]); 
    assign out[7152] = ~layer_0[9420]; 
    assign out[7153] = layer_0[974] ^ layer_0[6129]; 
    assign out[7154] = ~(layer_0[2601] ^ layer_0[10278]); 
    assign out[7155] = ~layer_0[6672] | (layer_0[6672] & layer_0[5327]); 
    assign out[7156] = ~(layer_0[10929] ^ layer_0[9171]); 
    assign out[7157] = layer_0[7275] ^ layer_0[6267]; 
    assign out[7158] = layer_0[778]; 
    assign out[7159] = ~layer_0[707]; 
    assign out[7160] = ~(layer_0[11629] ^ layer_0[10204]); 
    assign out[7161] = layer_0[5775] & ~layer_0[3822]; 
    assign out[7162] = ~(layer_0[11574] ^ layer_0[9871]); 
    assign out[7163] = ~layer_0[4244]; 
    assign out[7164] = layer_0[6325] ^ layer_0[5288]; 
    assign out[7165] = ~layer_0[4255]; 
    assign out[7166] = ~layer_0[10707] | (layer_0[10707] & layer_0[5595]); 
    assign out[7167] = ~(layer_0[8948] | layer_0[3239]); 
    assign out[7168] = layer_0[6474] | layer_0[6539]; 
    assign out[7169] = layer_0[8384]; 
    assign out[7170] = ~layer_0[3859] | (layer_0[8819] & layer_0[3859]); 
    assign out[7171] = layer_0[5766] & ~layer_0[5074]; 
    assign out[7172] = layer_0[7965] ^ layer_0[6143]; 
    assign out[7173] = ~layer_0[11879] | (layer_0[3563] & layer_0[11879]); 
    assign out[7174] = layer_0[301]; 
    assign out[7175] = ~(layer_0[5628] & layer_0[10677]); 
    assign out[7176] = ~(layer_0[8421] ^ layer_0[11327]); 
    assign out[7177] = layer_0[3378] ^ layer_0[3787]; 
    assign out[7178] = layer_0[3077] | layer_0[8505]; 
    assign out[7179] = ~(layer_0[1462] ^ layer_0[3463]); 
    assign out[7180] = ~(layer_0[10743] ^ layer_0[669]); 
    assign out[7181] = ~layer_0[5634] | (layer_0[5634] & layer_0[11172]); 
    assign out[7182] = ~(layer_0[406] & layer_0[1937]); 
    assign out[7183] = layer_0[8326]; 
    assign out[7184] = ~(layer_0[9104] ^ layer_0[11006]); 
    assign out[7185] = ~(layer_0[1136] & layer_0[6106]); 
    assign out[7186] = layer_0[11796]; 
    assign out[7187] = ~layer_0[5850] | (layer_0[5850] & layer_0[1834]); 
    assign out[7188] = ~(layer_0[7834] | layer_0[9693]); 
    assign out[7189] = ~layer_0[11543]; 
    assign out[7190] = layer_0[2923] | layer_0[7734]; 
    assign out[7191] = layer_0[10154] ^ layer_0[7561]; 
    assign out[7192] = layer_0[6541]; 
    assign out[7193] = layer_0[349] ^ layer_0[2613]; 
    assign out[7194] = layer_0[2655] | layer_0[2153]; 
    assign out[7195] = ~layer_0[2855] | (layer_0[2855] & layer_0[6837]); 
    assign out[7196] = ~(layer_0[89] ^ layer_0[3183]); 
    assign out[7197] = layer_0[10796]; 
    assign out[7198] = layer_0[4293] ^ layer_0[247]; 
    assign out[7199] = ~(layer_0[9978] ^ layer_0[9994]); 
    assign out[7200] = ~(layer_0[1400] ^ layer_0[11397]); 
    assign out[7201] = ~layer_0[3562]; 
    assign out[7202] = ~(layer_0[9260] ^ layer_0[2518]); 
    assign out[7203] = ~(layer_0[2542] & layer_0[7904]); 
    assign out[7204] = layer_0[8354] ^ layer_0[6032]; 
    assign out[7205] = ~(layer_0[6099] | layer_0[8105]); 
    assign out[7206] = layer_0[10895] ^ layer_0[6190]; 
    assign out[7207] = ~(layer_0[10509] | layer_0[1040]); 
    assign out[7208] = ~layer_0[1857]; 
    assign out[7209] = ~(layer_0[1920] ^ layer_0[5885]); 
    assign out[7210] = layer_0[9956]; 
    assign out[7211] = layer_0[8356] & ~layer_0[10093]; 
    assign out[7212] = layer_0[10949] & ~layer_0[6931]; 
    assign out[7213] = layer_0[15] & ~layer_0[11942]; 
    assign out[7214] = layer_0[3224]; 
    assign out[7215] = ~layer_0[5348]; 
    assign out[7216] = ~(layer_0[9457] | layer_0[8756]); 
    assign out[7217] = layer_0[11721]; 
    assign out[7218] = layer_0[901] & layer_0[10745]; 
    assign out[7219] = layer_0[11674]; 
    assign out[7220] = ~layer_0[7106]; 
    assign out[7221] = layer_0[11085] ^ layer_0[8105]; 
    assign out[7222] = ~layer_0[6096] | (layer_0[1048] & layer_0[6096]); 
    assign out[7223] = ~(layer_0[380] ^ layer_0[3806]); 
    assign out[7224] = layer_0[8770] ^ layer_0[11624]; 
    assign out[7225] = ~layer_0[6726]; 
    assign out[7226] = ~layer_0[8980] | (layer_0[8980] & layer_0[11969]); 
    assign out[7227] = ~layer_0[3652]; 
    assign out[7228] = layer_0[10995] & ~layer_0[3113]; 
    assign out[7229] = ~layer_0[4529]; 
    assign out[7230] = ~(layer_0[9408] ^ layer_0[8429]); 
    assign out[7231] = layer_0[11544]; 
    assign out[7232] = layer_0[627] ^ layer_0[7773]; 
    assign out[7233] = ~(layer_0[1926] ^ layer_0[3080]); 
    assign out[7234] = layer_0[6622] & ~layer_0[6603]; 
    assign out[7235] = ~(layer_0[257] ^ layer_0[9549]); 
    assign out[7236] = layer_0[1039] & ~layer_0[5684]; 
    assign out[7237] = layer_0[3747] ^ layer_0[1396]; 
    assign out[7238] = ~(layer_0[7785] | layer_0[6847]); 
    assign out[7239] = ~layer_0[8639] | (layer_0[2248] & layer_0[8639]); 
    assign out[7240] = layer_0[4006]; 
    assign out[7241] = layer_0[7008] ^ layer_0[8035]; 
    assign out[7242] = layer_0[4991] & layer_0[10510]; 
    assign out[7243] = layer_0[6271] & ~layer_0[11514]; 
    assign out[7244] = layer_0[7168] ^ layer_0[351]; 
    assign out[7245] = layer_0[11966] & ~layer_0[9757]; 
    assign out[7246] = ~(layer_0[9114] ^ layer_0[6784]); 
    assign out[7247] = layer_0[2729] ^ layer_0[9796]; 
    assign out[7248] = ~(layer_0[977] ^ layer_0[509]); 
    assign out[7249] = layer_0[10855] & ~layer_0[1403]; 
    assign out[7250] = ~(layer_0[11070] ^ layer_0[3484]); 
    assign out[7251] = layer_0[11728] & ~layer_0[2582]; 
    assign out[7252] = layer_0[9282] & ~layer_0[1793]; 
    assign out[7253] = ~(layer_0[4458] ^ layer_0[7305]); 
    assign out[7254] = layer_0[2139] ^ layer_0[2049]; 
    assign out[7255] = ~layer_0[5533]; 
    assign out[7256] = ~(layer_0[10400] ^ layer_0[2639]); 
    assign out[7257] = layer_0[782] ^ layer_0[3175]; 
    assign out[7258] = ~(layer_0[7663] ^ layer_0[4570]); 
    assign out[7259] = ~(layer_0[7028] | layer_0[7294]); 
    assign out[7260] = layer_0[4641]; 
    assign out[7261] = layer_0[2963] & ~layer_0[5969]; 
    assign out[7262] = ~(layer_0[5269] | layer_0[4358]); 
    assign out[7263] = layer_0[6083] & ~layer_0[9840]; 
    assign out[7264] = ~(layer_0[4625] ^ layer_0[8043]); 
    assign out[7265] = layer_0[9384] & ~layer_0[1317]; 
    assign out[7266] = ~(layer_0[7052] ^ layer_0[2619]); 
    assign out[7267] = layer_0[9658] ^ layer_0[5876]; 
    assign out[7268] = ~(layer_0[5122] ^ layer_0[937]); 
    assign out[7269] = layer_0[7379] & layer_0[8825]; 
    assign out[7270] = layer_0[9761] & layer_0[3593]; 
    assign out[7271] = ~(layer_0[8379] | layer_0[6426]); 
    assign out[7272] = layer_0[3075] ^ layer_0[9876]; 
    assign out[7273] = layer_0[9289] & layer_0[913]; 
    assign out[7274] = ~layer_0[2015]; 
    assign out[7275] = layer_0[6031] & ~layer_0[5037]; 
    assign out[7276] = layer_0[6227] ^ layer_0[4352]; 
    assign out[7277] = layer_0[9254] & layer_0[6710]; 
    assign out[7278] = layer_0[8231] ^ layer_0[2673]; 
    assign out[7279] = layer_0[9099]; 
    assign out[7280] = ~layer_0[1671]; 
    assign out[7281] = layer_0[4090] & ~layer_0[5100]; 
    assign out[7282] = ~(layer_0[11332] ^ layer_0[4167]); 
    assign out[7283] = ~(layer_0[5750] ^ layer_0[9882]); 
    assign out[7284] = layer_0[8088] & layer_0[2050]; 
    assign out[7285] = layer_0[303]; 
    assign out[7286] = ~(layer_0[10892] ^ layer_0[7084]); 
    assign out[7287] = layer_0[1782] ^ layer_0[1425]; 
    assign out[7288] = ~(layer_0[5372] ^ layer_0[875]); 
    assign out[7289] = ~(layer_0[7324] | layer_0[8316]); 
    assign out[7290] = layer_0[5205]; 
    assign out[7291] = layer_0[2939] ^ layer_0[6498]; 
    assign out[7292] = ~layer_0[6848] | (layer_0[6848] & layer_0[8069]); 
    assign out[7293] = layer_0[9040] & ~layer_0[7542]; 
    assign out[7294] = layer_0[921] | layer_0[6690]; 
    assign out[7295] = ~(layer_0[2026] ^ layer_0[8996]); 
    assign out[7296] = ~(layer_0[8007] | layer_0[9447]); 
    assign out[7297] = ~layer_0[9844] | (layer_0[3104] & layer_0[9844]); 
    assign out[7298] = ~(layer_0[5235] ^ layer_0[10984]); 
    assign out[7299] = ~layer_0[3876]; 
    assign out[7300] = layer_0[5177] & ~layer_0[3356]; 
    assign out[7301] = layer_0[4048] ^ layer_0[6139]; 
    assign out[7302] = ~layer_0[3171]; 
    assign out[7303] = ~(layer_0[2308] | layer_0[4141]); 
    assign out[7304] = ~(layer_0[4249] ^ layer_0[1316]); 
    assign out[7305] = ~(layer_0[3278] ^ layer_0[4694]); 
    assign out[7306] = ~layer_0[5884] | (layer_0[5884] & layer_0[10369]); 
    assign out[7307] = layer_0[10414]; 
    assign out[7308] = layer_0[5060] ^ layer_0[9801]; 
    assign out[7309] = ~layer_0[7583]; 
    assign out[7310] = ~(layer_0[6834] & layer_0[3383]); 
    assign out[7311] = ~(layer_0[4089] ^ layer_0[8814]); 
    assign out[7312] = ~layer_0[11656]; 
    assign out[7313] = ~layer_0[10913]; 
    assign out[7314] = ~(layer_0[1651] | layer_0[5904]); 
    assign out[7315] = layer_0[11793] ^ layer_0[10025]; 
    assign out[7316] = layer_0[8602] ^ layer_0[11588]; 
    assign out[7317] = layer_0[4805] & ~layer_0[1505]; 
    assign out[7318] = layer_0[3550] & ~layer_0[6933]; 
    assign out[7319] = layer_0[557] & ~layer_0[9881]; 
    assign out[7320] = layer_0[7338] & layer_0[9787]; 
    assign out[7321] = layer_0[265] ^ layer_0[5117]; 
    assign out[7322] = layer_0[7907] & layer_0[10830]; 
    assign out[7323] = ~(layer_0[6157] | layer_0[1101]); 
    assign out[7324] = ~(layer_0[11772] | layer_0[7608]); 
    assign out[7325] = layer_0[6289] & layer_0[11441]; 
    assign out[7326] = layer_0[5393] & layer_0[10861]; 
    assign out[7327] = layer_0[8633] ^ layer_0[6828]; 
    assign out[7328] = layer_0[7915] ^ layer_0[3686]; 
    assign out[7329] = ~(layer_0[9178] ^ layer_0[2108]); 
    assign out[7330] = layer_0[1624] ^ layer_0[11751]; 
    assign out[7331] = ~(layer_0[8448] | layer_0[7659]); 
    assign out[7332] = layer_0[9666] & ~layer_0[11271]; 
    assign out[7333] = ~layer_0[4733]; 
    assign out[7334] = layer_0[11635] & ~layer_0[506]; 
    assign out[7335] = layer_0[4569] | layer_0[2850]; 
    assign out[7336] = layer_0[3280] & layer_0[7002]; 
    assign out[7337] = ~layer_0[4095]; 
    assign out[7338] = ~layer_0[2982]; 
    assign out[7339] = ~(layer_0[8841] ^ layer_0[5169]); 
    assign out[7340] = ~(layer_0[8853] ^ layer_0[9229]); 
    assign out[7341] = ~(layer_0[1704] ^ layer_0[10809]); 
    assign out[7342] = ~layer_0[10496]; 
    assign out[7343] = layer_0[8376] ^ layer_0[5428]; 
    assign out[7344] = layer_0[1463] ^ layer_0[11770]; 
    assign out[7345] = ~(layer_0[8764] | layer_0[1778]); 
    assign out[7346] = layer_0[7649] & ~layer_0[11783]; 
    assign out[7347] = layer_0[1051] ^ layer_0[3852]; 
    assign out[7348] = layer_0[5116] & ~layer_0[4798]; 
    assign out[7349] = layer_0[140] & ~layer_0[5413]; 
    assign out[7350] = ~layer_0[1410]; 
    assign out[7351] = ~(layer_0[318] ^ layer_0[11579]); 
    assign out[7352] = layer_0[9237] & layer_0[2316]; 
    assign out[7353] = ~(layer_0[1362] & layer_0[8437]); 
    assign out[7354] = ~(layer_0[5074] ^ layer_0[3229]); 
    assign out[7355] = layer_0[4586] & layer_0[4954]; 
    assign out[7356] = ~(layer_0[6026] ^ layer_0[11839]); 
    assign out[7357] = ~layer_0[2123]; 
    assign out[7358] = layer_0[8580] ^ layer_0[10860]; 
    assign out[7359] = layer_0[4432] & layer_0[7019]; 
    assign out[7360] = layer_0[1860] ^ layer_0[8953]; 
    assign out[7361] = ~(layer_0[7689] ^ layer_0[9527]); 
    assign out[7362] = layer_0[5335] ^ layer_0[5295]; 
    assign out[7363] = layer_0[5158] ^ layer_0[3526]; 
    assign out[7364] = ~(layer_0[9679] ^ layer_0[6876]); 
    assign out[7365] = ~(layer_0[918] | layer_0[3204]); 
    assign out[7366] = layer_0[2073] ^ layer_0[4452]; 
    assign out[7367] = ~(layer_0[10637] ^ layer_0[7491]); 
    assign out[7368] = ~(layer_0[510] | layer_0[7004]); 
    assign out[7369] = layer_0[4666] ^ layer_0[7594]; 
    assign out[7370] = ~(layer_0[7330] ^ layer_0[3009]); 
    assign out[7371] = layer_0[33] ^ layer_0[11129]; 
    assign out[7372] = ~layer_0[9622]; 
    assign out[7373] = ~(layer_0[9719] & layer_0[3574]); 
    assign out[7374] = layer_0[569] & ~layer_0[4446]; 
    assign out[7375] = ~layer_0[10916]; 
    assign out[7376] = layer_0[7448] ^ layer_0[9858]; 
    assign out[7377] = layer_0[432] & ~layer_0[7117]; 
    assign out[7378] = layer_0[2210] | layer_0[2802]; 
    assign out[7379] = ~(layer_0[1191] ^ layer_0[2430]); 
    assign out[7380] = layer_0[4432] & ~layer_0[11411]; 
    assign out[7381] = layer_0[3606] & layer_0[3458]; 
    assign out[7382] = layer_0[2131] ^ layer_0[10018]; 
    assign out[7383] = ~(layer_0[6751] | layer_0[5797]); 
    assign out[7384] = layer_0[3551] & ~layer_0[7220]; 
    assign out[7385] = ~(layer_0[7692] ^ layer_0[7377]); 
    assign out[7386] = ~layer_0[9841]; 
    assign out[7387] = ~(layer_0[9018] ^ layer_0[6889]); 
    assign out[7388] = layer_0[433] ^ layer_0[3765]; 
    assign out[7389] = ~layer_0[6203]; 
    assign out[7390] = ~layer_0[9920]; 
    assign out[7391] = layer_0[11258] & ~layer_0[10016]; 
    assign out[7392] = layer_0[3142] & layer_0[8930]; 
    assign out[7393] = layer_0[9017] ^ layer_0[2437]; 
    assign out[7394] = ~layer_0[2124]; 
    assign out[7395] = layer_0[1736] & ~layer_0[9307]; 
    assign out[7396] = layer_0[6789]; 
    assign out[7397] = ~(layer_0[3708] ^ layer_0[6194]); 
    assign out[7398] = layer_0[4204] & layer_0[592]; 
    assign out[7399] = layer_0[7315] ^ layer_0[6517]; 
    assign out[7400] = ~layer_0[7353]; 
    assign out[7401] = layer_0[5338] & ~layer_0[5648]; 
    assign out[7402] = layer_0[6007] ^ layer_0[2329]; 
    assign out[7403] = ~layer_0[6272]; 
    assign out[7404] = ~(layer_0[4300] ^ layer_0[3835]); 
    assign out[7405] = layer_0[2162] ^ layer_0[10250]; 
    assign out[7406] = layer_0[11227] ^ layer_0[9125]; 
    assign out[7407] = ~(layer_0[9187] ^ layer_0[4908]); 
    assign out[7408] = layer_0[8409] ^ layer_0[4215]; 
    assign out[7409] = layer_0[9459] ^ layer_0[7624]; 
    assign out[7410] = layer_0[8060] & ~layer_0[119]; 
    assign out[7411] = ~(layer_0[11974] ^ layer_0[8317]); 
    assign out[7412] = layer_0[7805] & ~layer_0[5859]; 
    assign out[7413] = layer_0[6929] & ~layer_0[2068]; 
    assign out[7414] = layer_0[9995] ^ layer_0[5197]; 
    assign out[7415] = layer_0[7961] & layer_0[7261]; 
    assign out[7416] = ~(layer_0[11571] ^ layer_0[7249]); 
    assign out[7417] = layer_0[9716] & ~layer_0[1749]; 
    assign out[7418] = layer_0[5307] ^ layer_0[1824]; 
    assign out[7419] = ~layer_0[2376] | (layer_0[2376] & layer_0[9768]); 
    assign out[7420] = ~(layer_0[9975] | layer_0[9312]); 
    assign out[7421] = ~layer_0[8063]; 
    assign out[7422] = ~(layer_0[10405] | layer_0[10951]); 
    assign out[7423] = ~(layer_0[5870] ^ layer_0[3294]); 
    assign out[7424] = layer_0[10617] ^ layer_0[3729]; 
    assign out[7425] = ~(layer_0[3823] ^ layer_0[2025]); 
    assign out[7426] = layer_0[8708] & ~layer_0[10258]; 
    assign out[7427] = layer_0[113]; 
    assign out[7428] = layer_0[5342] ^ layer_0[4280]; 
    assign out[7429] = layer_0[8416] & ~layer_0[5047]; 
    assign out[7430] = ~(layer_0[2168] & layer_0[41]); 
    assign out[7431] = ~(layer_0[2448] ^ layer_0[1820]); 
    assign out[7432] = layer_0[2994] & layer_0[3101]; 
    assign out[7433] = layer_0[9028]; 
    assign out[7434] = layer_0[7843] ^ layer_0[5854]; 
    assign out[7435] = ~(layer_0[4951] ^ layer_0[2739]); 
    assign out[7436] = ~(layer_0[6011] ^ layer_0[11594]); 
    assign out[7437] = layer_0[7524]; 
    assign out[7438] = layer_0[8412]; 
    assign out[7439] = ~layer_0[10630]; 
    assign out[7440] = ~layer_0[5437]; 
    assign out[7441] = layer_0[3316] & ~layer_0[1776]; 
    assign out[7442] = ~(layer_0[3503] | layer_0[844]); 
    assign out[7443] = layer_0[8332] & ~layer_0[8097]; 
    assign out[7444] = layer_0[9493]; 
    assign out[7445] = layer_0[5245] & ~layer_0[1254]; 
    assign out[7446] = layer_0[9646] & ~layer_0[5679]; 
    assign out[7447] = ~layer_0[7412] | (layer_0[3393] & layer_0[7412]); 
    assign out[7448] = layer_0[9750]; 
    assign out[7449] = layer_0[9210] & layer_0[5419]; 
    assign out[7450] = layer_0[4774] & ~layer_0[3521]; 
    assign out[7451] = layer_0[4294] & layer_0[9446]; 
    assign out[7452] = layer_0[4102]; 
    assign out[7453] = layer_0[7512] ^ layer_0[7732]; 
    assign out[7454] = ~(layer_0[2682] | layer_0[1881]); 
    assign out[7455] = ~layer_0[6544]; 
    assign out[7456] = ~(layer_0[2398] ^ layer_0[9362]); 
    assign out[7457] = layer_0[4004] & ~layer_0[7892]; 
    assign out[7458] = ~(layer_0[5902] ^ layer_0[7560]); 
    assign out[7459] = ~(layer_0[2426] | layer_0[8530]); 
    assign out[7460] = layer_0[8304] ^ layer_0[1908]; 
    assign out[7461] = ~(layer_0[773] | layer_0[2617]); 
    assign out[7462] = ~(layer_0[10179] ^ layer_0[10609]); 
    assign out[7463] = ~(layer_0[1638] & layer_0[3088]); 
    assign out[7464] = ~layer_0[8876] | (layer_0[453] & layer_0[8876]); 
    assign out[7465] = layer_0[8583] ^ layer_0[2257]; 
    assign out[7466] = layer_0[10236] ^ layer_0[10823]; 
    assign out[7467] = ~layer_0[10146]; 
    assign out[7468] = ~(layer_0[7611] ^ layer_0[6998]); 
    assign out[7469] = layer_0[4099] ^ layer_0[10242]; 
    assign out[7470] = ~(layer_0[7458] ^ layer_0[3933]); 
    assign out[7471] = ~layer_0[7782]; 
    assign out[7472] = layer_0[9094] & layer_0[5793]; 
    assign out[7473] = ~(layer_0[443] | layer_0[1268]); 
    assign out[7474] = layer_0[5183] ^ layer_0[11283]; 
    assign out[7475] = layer_0[11638] ^ layer_0[1406]; 
    assign out[7476] = layer_0[3175] & ~layer_0[6137]; 
    assign out[7477] = ~(layer_0[6392] ^ layer_0[11733]); 
    assign out[7478] = layer_0[1549] & ~layer_0[6645]; 
    assign out[7479] = layer_0[9205] & layer_0[1469]; 
    assign out[7480] = ~(layer_0[360] | layer_0[10593]); 
    assign out[7481] = ~layer_0[4401]; 
    assign out[7482] = layer_0[9445] & ~layer_0[11628]; 
    assign out[7483] = layer_0[3696] ^ layer_0[795]; 
    assign out[7484] = ~(layer_0[11260] | layer_0[4160]); 
    assign out[7485] = ~(layer_0[3567] ^ layer_0[7657]); 
    assign out[7486] = layer_0[3514]; 
    assign out[7487] = layer_0[331] ^ layer_0[3962]; 
    assign out[7488] = ~(layer_0[10150] ^ layer_0[5130]); 
    assign out[7489] = layer_0[10635] & ~layer_0[10193]; 
    assign out[7490] = layer_0[2547] & ~layer_0[3589]; 
    assign out[7491] = ~layer_0[4867]; 
    assign out[7492] = ~layer_0[8139]; 
    assign out[7493] = layer_0[5528] ^ layer_0[9195]; 
    assign out[7494] = layer_0[6757] & layer_0[808]; 
    assign out[7495] = ~(layer_0[340] | layer_0[7848]); 
    assign out[7496] = layer_0[11348] & layer_0[7330]; 
    assign out[7497] = ~(layer_0[4779] | layer_0[9134]); 
    assign out[7498] = layer_0[4346] & layer_0[10828]; 
    assign out[7499] = ~(layer_0[3306] ^ layer_0[8822]); 
    assign out[7500] = layer_0[6486] ^ layer_0[10583]; 
    assign out[7501] = ~layer_0[6302]; 
    assign out[7502] = layer_0[3255] & ~layer_0[7427]; 
    assign out[7503] = layer_0[11113]; 
    assign out[7504] = ~layer_0[5377] | (layer_0[5936] & layer_0[5377]); 
    assign out[7505] = layer_0[7972] & ~layer_0[9432]; 
    assign out[7506] = ~layer_0[8303]; 
    assign out[7507] = ~(layer_0[6778] ^ layer_0[8355]); 
    assign out[7508] = layer_0[7834] ^ layer_0[1766]; 
    assign out[7509] = layer_0[1676] ^ layer_0[172]; 
    assign out[7510] = layer_0[3641] ^ layer_0[5123]; 
    assign out[7511] = layer_0[4327]; 
    assign out[7512] = layer_0[982]; 
    assign out[7513] = layer_0[11969] | layer_0[6819]; 
    assign out[7514] = ~layer_0[1524] | (layer_0[5720] & layer_0[1524]); 
    assign out[7515] = layer_0[10474] & layer_0[11743]; 
    assign out[7516] = layer_0[11696] ^ layer_0[4979]; 
    assign out[7517] = ~(layer_0[7187] | layer_0[11142]); 
    assign out[7518] = layer_0[9235] & layer_0[84]; 
    assign out[7519] = layer_0[9531] ^ layer_0[9741]; 
    assign out[7520] = ~(layer_0[10789] | layer_0[10764]); 
    assign out[7521] = ~(layer_0[7918] | layer_0[10294]); 
    assign out[7522] = ~(layer_0[5748] ^ layer_0[2788]); 
    assign out[7523] = layer_0[3849] & layer_0[3002]; 
    assign out[7524] = ~layer_0[1602] | (layer_0[8386] & layer_0[1602]); 
    assign out[7525] = ~layer_0[4392]; 
    assign out[7526] = layer_0[5035] ^ layer_0[5631]; 
    assign out[7527] = ~(layer_0[488] ^ layer_0[11593]); 
    assign out[7528] = layer_0[3231]; 
    assign out[7529] = ~layer_0[556]; 
    assign out[7530] = ~(layer_0[1634] ^ layer_0[3525]); 
    assign out[7531] = layer_0[5265] & ~layer_0[4480]; 
    assign out[7532] = layer_0[6141] ^ layer_0[4186]; 
    assign out[7533] = ~layer_0[11955]; 
    assign out[7534] = ~(layer_0[3031] ^ layer_0[2675]); 
    assign out[7535] = ~(layer_0[10758] ^ layer_0[10607]); 
    assign out[7536] = layer_0[11483]; 
    assign out[7537] = layer_0[8255] ^ layer_0[9714]; 
    assign out[7538] = layer_0[7306] | layer_0[7196]; 
    assign out[7539] = layer_0[9398]; 
    assign out[7540] = layer_0[9142] ^ layer_0[1870]; 
    assign out[7541] = layer_0[8630] & layer_0[7735]; 
    assign out[7542] = ~layer_0[11566]; 
    assign out[7543] = layer_0[4585] ^ layer_0[6248]; 
    assign out[7544] = ~(layer_0[5349] ^ layer_0[1141]); 
    assign out[7545] = layer_0[7529] | layer_0[5882]; 
    assign out[7546] = layer_0[3203] & ~layer_0[11216]; 
    assign out[7547] = layer_0[5249]; 
    assign out[7548] = ~layer_0[3455]; 
    assign out[7549] = layer_0[8411] & ~layer_0[8888]; 
    assign out[7550] = ~(layer_0[11063] ^ layer_0[1484]); 
    assign out[7551] = ~(layer_0[9980] ^ layer_0[6178]); 
    assign out[7552] = layer_0[7800] ^ layer_0[4117]; 
    assign out[7553] = layer_0[7775] & ~layer_0[3432]; 
    assign out[7554] = ~layer_0[457] | (layer_0[457] & layer_0[5550]); 
    assign out[7555] = layer_0[4533] & ~layer_0[820]; 
    assign out[7556] = layer_0[2156] ^ layer_0[8027]; 
    assign out[7557] = ~(layer_0[2382] & layer_0[3361]); 
    assign out[7558] = layer_0[3507] ^ layer_0[939]; 
    assign out[7559] = layer_0[11837]; 
    assign out[7560] = ~(layer_0[9368] ^ layer_0[4974]); 
    assign out[7561] = ~(layer_0[3648] | layer_0[1540]); 
    assign out[7562] = ~layer_0[9179] | (layer_0[3812] & layer_0[9179]); 
    assign out[7563] = layer_0[9933] ^ layer_0[3827]; 
    assign out[7564] = layer_0[2905] ^ layer_0[9620]; 
    assign out[7565] = layer_0[7646] & ~layer_0[3819]; 
    assign out[7566] = ~(layer_0[8536] | layer_0[6776]); 
    assign out[7567] = ~(layer_0[7421] ^ layer_0[1843]); 
    assign out[7568] = ~(layer_0[5104] | layer_0[1059]); 
    assign out[7569] = ~layer_0[5454]; 
    assign out[7570] = layer_0[5093] & ~layer_0[195]; 
    assign out[7571] = layer_0[6417] ^ layer_0[9912]; 
    assign out[7572] = layer_0[8845] ^ layer_0[4765]; 
    assign out[7573] = layer_0[507]; 
    assign out[7574] = layer_0[10654] & ~layer_0[8911]; 
    assign out[7575] = layer_0[5173] & ~layer_0[7600]; 
    assign out[7576] = ~(layer_0[8244] | layer_0[9816]); 
    assign out[7577] = ~layer_0[6715]; 
    assign out[7578] = layer_0[10158]; 
    assign out[7579] = ~(layer_0[10844] ^ layer_0[6942]); 
    assign out[7580] = ~(layer_0[10433] & layer_0[3439]); 
    assign out[7581] = ~(layer_0[7607] ^ layer_0[7003]); 
    assign out[7582] = ~layer_0[11850]; 
    assign out[7583] = layer_0[4661] & layer_0[9068]; 
    assign out[7584] = layer_0[11692]; 
    assign out[7585] = layer_0[8044]; 
    assign out[7586] = ~(layer_0[11905] | layer_0[1839]); 
    assign out[7587] = ~(layer_0[11511] ^ layer_0[3309]); 
    assign out[7588] = 1'b0; 
    assign out[7589] = ~(layer_0[4018] ^ layer_0[3529]); 
    assign out[7590] = layer_0[3082] & ~layer_0[8662]; 
    assign out[7591] = ~(layer_0[8115] | layer_0[4782]); 
    assign out[7592] = ~(layer_0[9642] | layer_0[9441]); 
    assign out[7593] = ~layer_0[1382]; 
    assign out[7594] = layer_0[1700] & ~layer_0[6232]; 
    assign out[7595] = layer_0[6069] ^ layer_0[6610]; 
    assign out[7596] = ~layer_0[8070] | (layer_0[1230] & layer_0[8070]); 
    assign out[7597] = ~(layer_0[3527] | layer_0[10760]); 
    assign out[7598] = ~(layer_0[1659] ^ layer_0[9151]); 
    assign out[7599] = layer_0[7067] ^ layer_0[3493]; 
    assign out[7600] = ~(layer_0[1336] ^ layer_0[10556]); 
    assign out[7601] = layer_0[7435] & ~layer_0[4986]; 
    assign out[7602] = layer_0[9764]; 
    assign out[7603] = ~(layer_0[195] | layer_0[5229]); 
    assign out[7604] = layer_0[11343] & ~layer_0[6261]; 
    assign out[7605] = layer_0[6479]; 
    assign out[7606] = layer_0[5467] ^ layer_0[40]; 
    assign out[7607] = layer_0[5632]; 
    assign out[7608] = layer_0[311] ^ layer_0[2933]; 
    assign out[7609] = layer_0[1019] ^ layer_0[11121]; 
    assign out[7610] = layer_0[1454]; 
    assign out[7611] = 1'b1; 
    assign out[7612] = layer_0[5490] & ~layer_0[3065]; 
    assign out[7613] = layer_0[11507]; 
    assign out[7614] = ~layer_0[1422] | (layer_0[6222] & layer_0[1422]); 
    assign out[7615] = ~(layer_0[3465] ^ layer_0[10837]); 
    assign out[7616] = layer_0[9155] ^ layer_0[7231]; 
    assign out[7617] = ~(layer_0[7061] | layer_0[1595]); 
    assign out[7618] = ~layer_0[148] | (layer_0[148] & layer_0[8055]); 
    assign out[7619] = ~(layer_0[7316] ^ layer_0[8264]); 
    assign out[7620] = layer_0[5196] & ~layer_0[9749]; 
    assign out[7621] = layer_0[10736] & ~layer_0[7683]; 
    assign out[7622] = layer_0[631] ^ layer_0[5597]; 
    assign out[7623] = layer_0[9907] & ~layer_0[11132]; 
    assign out[7624] = ~(layer_0[616] | layer_0[1603]); 
    assign out[7625] = layer_0[11201] & layer_0[9778]; 
    assign out[7626] = layer_0[11503] & layer_0[5958]; 
    assign out[7627] = ~layer_0[5535] | (layer_0[5535] & layer_0[10919]); 
    assign out[7628] = ~(layer_0[11938] ^ layer_0[7038]); 
    assign out[7629] = layer_0[7637] & ~layer_0[1040]; 
    assign out[7630] = layer_0[678] & ~layer_0[11494]; 
    assign out[7631] = layer_0[6160] & layer_0[6234]; 
    assign out[7632] = ~(layer_0[9020] | layer_0[9715]); 
    assign out[7633] = layer_0[3739] & ~layer_0[3412]; 
    assign out[7634] = ~layer_0[1895]; 
    assign out[7635] = layer_0[203] & layer_0[1981]; 
    assign out[7636] = layer_0[4649] ^ layer_0[2978]; 
    assign out[7637] = layer_0[11764]; 
    assign out[7638] = layer_0[4202] ^ layer_0[6356]; 
    assign out[7639] = layer_0[8579]; 
    assign out[7640] = ~(layer_0[6475] ^ layer_0[11665]); 
    assign out[7641] = layer_0[1805] & ~layer_0[7488]; 
    assign out[7642] = layer_0[11095] & layer_0[2742]; 
    assign out[7643] = layer_0[10874] & layer_0[202]; 
    assign out[7644] = layer_0[3468] & ~layer_0[4727]; 
    assign out[7645] = ~(layer_0[8344] ^ layer_0[10760]); 
    assign out[7646] = ~layer_0[7804]; 
    assign out[7647] = layer_0[7113] & layer_0[8660]; 
    assign out[7648] = layer_0[2562] ^ layer_0[9088]; 
    assign out[7649] = layer_0[1107] & ~layer_0[1535]; 
    assign out[7650] = layer_0[9441] & layer_0[4341]; 
    assign out[7651] = ~(layer_0[4821] ^ layer_0[6771]); 
    assign out[7652] = ~layer_0[10168] | (layer_0[4588] & layer_0[10168]); 
    assign out[7653] = ~(layer_0[4069] ^ layer_0[7801]); 
    assign out[7654] = ~(layer_0[3076] | layer_0[5899]); 
    assign out[7655] = ~(layer_0[516] ^ layer_0[9556]); 
    assign out[7656] = layer_0[9821] ^ layer_0[3325]; 
    assign out[7657] = layer_0[1772] ^ layer_0[1483]; 
    assign out[7658] = layer_0[3267] & ~layer_0[10020]; 
    assign out[7659] = layer_0[10989] & layer_0[10463]; 
    assign out[7660] = ~(layer_0[9653] | layer_0[10902]); 
    assign out[7661] = layer_0[4553] & layer_0[1332]; 
    assign out[7662] = layer_0[6543] ^ layer_0[11371]; 
    assign out[7663] = layer_0[2808] & layer_0[10490]; 
    assign out[7664] = layer_0[10328] ^ layer_0[7399]; 
    assign out[7665] = ~(layer_0[2900] | layer_0[4503]); 
    assign out[7666] = layer_0[11607] ^ layer_0[9822]; 
    assign out[7667] = layer_0[5751] | layer_0[4990]; 
    assign out[7668] = layer_0[222] & ~layer_0[5096]; 
    assign out[7669] = layer_0[4713] & ~layer_0[8845]; 
    assign out[7670] = layer_0[8394] ^ layer_0[7712]; 
    assign out[7671] = layer_0[7370] ^ layer_0[1002]; 
    assign out[7672] = ~(layer_0[3402] ^ layer_0[10221]); 
    assign out[7673] = ~(layer_0[6947] ^ layer_0[8548]); 
    assign out[7674] = layer_0[8265] & ~layer_0[8712]; 
    assign out[7675] = layer_0[2647] | layer_0[7006]; 
    assign out[7676] = layer_0[4790] ^ layer_0[1786]; 
    assign out[7677] = layer_0[3857] & layer_0[6369]; 
    assign out[7678] = layer_0[5536]; 
    assign out[7679] = ~(layer_0[1878] & layer_0[7852]); 
    assign out[7680] = ~layer_0[9333]; 
    assign out[7681] = layer_0[3392] & layer_0[1069]; 
    assign out[7682] = layer_0[6450] ^ layer_0[847]; 
    assign out[7683] = ~(layer_0[2925] | layer_0[492]); 
    assign out[7684] = layer_0[7354] & layer_0[7269]; 
    assign out[7685] = layer_0[4002] ^ layer_0[965]; 
    assign out[7686] = layer_0[4236] & ~layer_0[1129]; 
    assign out[7687] = layer_0[2888] & ~layer_0[10217]; 
    assign out[7688] = layer_0[4913] ^ layer_0[3670]; 
    assign out[7689] = ~(layer_0[2122] & layer_0[2515]); 
    assign out[7690] = ~(layer_0[5056] ^ layer_0[7233]); 
    assign out[7691] = layer_0[7798]; 
    assign out[7692] = layer_0[5389] & layer_0[3988]; 
    assign out[7693] = layer_0[1539] & ~layer_0[362]; 
    assign out[7694] = layer_0[7080] & layer_0[8493]; 
    assign out[7695] = layer_0[3913] & layer_0[5726]; 
    assign out[7696] = layer_0[2403] ^ layer_0[8588]; 
    assign out[7697] = ~(layer_0[3469] ^ layer_0[5048]); 
    assign out[7698] = layer_0[3377] & layer_0[11193]; 
    assign out[7699] = ~(layer_0[670] ^ layer_0[6971]); 
    assign out[7700] = layer_0[4706] ^ layer_0[4057]; 
    assign out[7701] = layer_0[6755] ^ layer_0[8305]; 
    assign out[7702] = layer_0[8541] & layer_0[7714]; 
    assign out[7703] = layer_0[5515] & layer_0[3014]; 
    assign out[7704] = ~(layer_0[126] ^ layer_0[522]); 
    assign out[7705] = layer_0[11794] & layer_0[1593]; 
    assign out[7706] = layer_0[11833]; 
    assign out[7707] = layer_0[2741] & ~layer_0[6077]; 
    assign out[7708] = layer_0[8931] | layer_0[1534]; 
    assign out[7709] = layer_0[8826]; 
    assign out[7710] = layer_0[2160]; 
    assign out[7711] = ~(layer_0[831] | layer_0[10570]); 
    assign out[7712] = ~(layer_0[11172] | layer_0[7147]); 
    assign out[7713] = layer_0[4624] & layer_0[968]; 
    assign out[7714] = layer_0[6983] & layer_0[3280]; 
    assign out[7715] = ~(layer_0[11771] | layer_0[11667]); 
    assign out[7716] = ~(layer_0[2896] | layer_0[8390]); 
    assign out[7717] = ~layer_0[10578]; 
    assign out[7718] = layer_0[5706] & ~layer_0[10765]; 
    assign out[7719] = layer_0[10522] & ~layer_0[10067]; 
    assign out[7720] = layer_0[11928] ^ layer_0[7971]; 
    assign out[7721] = layer_0[11123] ^ layer_0[10669]; 
    assign out[7722] = ~layer_0[9219]; 
    assign out[7723] = ~(layer_0[8522] | layer_0[7525]); 
    assign out[7724] = ~(layer_0[10953] ^ layer_0[4859]); 
    assign out[7725] = layer_0[4965]; 
    assign out[7726] = ~(layer_0[4319] ^ layer_0[3268]); 
    assign out[7727] = ~(layer_0[6292] & layer_0[3357]); 
    assign out[7728] = layer_0[6984] & ~layer_0[9628]; 
    assign out[7729] = ~(layer_0[4324] | layer_0[4693]); 
    assign out[7730] = layer_0[641] ^ layer_0[8943]; 
    assign out[7731] = layer_0[417]; 
    assign out[7732] = ~(layer_0[3009] ^ layer_0[431]); 
    assign out[7733] = layer_0[1139] | layer_0[10827]; 
    assign out[7734] = ~layer_0[1308]; 
    assign out[7735] = layer_0[2401]; 
    assign out[7736] = layer_0[7180] & ~layer_0[1728]; 
    assign out[7737] = layer_0[6690] & layer_0[7344]; 
    assign out[7738] = layer_0[5617] ^ layer_0[5786]; 
    assign out[7739] = layer_0[6903] & ~layer_0[9846]; 
    assign out[7740] = layer_0[8434] & ~layer_0[5742]; 
    assign out[7741] = layer_0[2708] & layer_0[11034]; 
    assign out[7742] = ~(layer_0[9463] ^ layer_0[11002]); 
    assign out[7743] = ~layer_0[7429]; 
    assign out[7744] = ~(layer_0[11343] ^ layer_0[7650]); 
    assign out[7745] = layer_0[9363] & ~layer_0[3846]; 
    assign out[7746] = ~(layer_0[4138] ^ layer_0[9332]); 
    assign out[7747] = layer_0[405] ^ layer_0[8197]; 
    assign out[7748] = layer_0[9964] & ~layer_0[4874]; 
    assign out[7749] = ~(layer_0[11449] | layer_0[11386]); 
    assign out[7750] = ~layer_0[1948]; 
    assign out[7751] = layer_0[9870]; 
    assign out[7752] = ~(layer_0[2330] | layer_0[1840]); 
    assign out[7753] = layer_0[5421]; 
    assign out[7754] = layer_0[4466] ^ layer_0[9067]; 
    assign out[7755] = layer_0[7048] & ~layer_0[3478]; 
    assign out[7756] = layer_0[5450] ^ layer_0[6545]; 
    assign out[7757] = ~(layer_0[7392] | layer_0[8245]); 
    assign out[7758] = layer_0[5971] ^ layer_0[3253]; 
    assign out[7759] = ~layer_0[10912]; 
    assign out[7760] = layer_0[4029] & ~layer_0[3806]; 
    assign out[7761] = ~(layer_0[6330] | layer_0[5530]); 
    assign out[7762] = layer_0[9640]; 
    assign out[7763] = layer_0[8166] & ~layer_0[5878]; 
    assign out[7764] = layer_0[3900] ^ layer_0[6485]; 
    assign out[7765] = ~(layer_0[2063] & layer_0[10074]); 
    assign out[7766] = ~(layer_0[7409] ^ layer_0[4503]); 
    assign out[7767] = layer_0[165]; 
    assign out[7768] = ~layer_0[11166]; 
    assign out[7769] = ~(layer_0[7779] ^ layer_0[6125]); 
    assign out[7770] = layer_0[4949] ^ layer_0[7334]; 
    assign out[7771] = ~(layer_0[1412] | layer_0[1943]); 
    assign out[7772] = ~(layer_0[2640] ^ layer_0[10640]); 
    assign out[7773] = layer_0[8223] ^ layer_0[11744]; 
    assign out[7774] = ~(layer_0[799] ^ layer_0[9176]); 
    assign out[7775] = ~layer_0[1672] | (layer_0[1672] & layer_0[2769]); 
    assign out[7776] = ~(layer_0[7341] ^ layer_0[9934]); 
    assign out[7777] = 1'b0; 
    assign out[7778] = layer_0[6866]; 
    assign out[7779] = layer_0[3969]; 
    assign out[7780] = ~layer_0[8764]; 
    assign out[7781] = layer_0[11977] & ~layer_0[9112]; 
    assign out[7782] = layer_0[9931] & ~layer_0[9348]; 
    assign out[7783] = ~(layer_0[1063] ^ layer_0[9686]); 
    assign out[7784] = layer_0[1663] & layer_0[5520]; 
    assign out[7785] = layer_0[4102] & ~layer_0[4337]; 
    assign out[7786] = ~(layer_0[1126] ^ layer_0[10662]); 
    assign out[7787] = ~(layer_0[2339] ^ layer_0[7970]); 
    assign out[7788] = ~(layer_0[6552] ^ layer_0[9387]); 
    assign out[7789] = layer_0[11355] ^ layer_0[10933]; 
    assign out[7790] = layer_0[7301]; 
    assign out[7791] = ~(layer_0[4890] ^ layer_0[1238]); 
    assign out[7792] = ~(layer_0[2086] ^ layer_0[8415]); 
    assign out[7793] = layer_0[3775] ^ layer_0[4119]; 
    assign out[7794] = layer_0[7300] & ~layer_0[11413]; 
    assign out[7795] = ~(layer_0[282] ^ layer_0[7214]); 
    assign out[7796] = ~(layer_0[660] ^ layer_0[9413]); 
    assign out[7797] = layer_0[8342]; 
    assign out[7798] = layer_0[3539]; 
    assign out[7799] = ~(layer_0[10336] ^ layer_0[5979]); 
    assign out[7800] = layer_0[6826] & ~layer_0[11378]; 
    assign out[7801] = ~layer_0[7091]; 
    assign out[7802] = layer_0[5778] ^ layer_0[781]; 
    assign out[7803] = layer_0[1569] & ~layer_0[9687]; 
    assign out[7804] = layer_0[9733] ^ layer_0[5735]; 
    assign out[7805] = ~(layer_0[579] | layer_0[3260]); 
    assign out[7806] = layer_0[2539] ^ layer_0[2424]; 
    assign out[7807] = layer_0[3815] | layer_0[11825]; 
    assign out[7808] = layer_0[304] & ~layer_0[4817]; 
    assign out[7809] = layer_0[6336]; 
    assign out[7810] = ~(layer_0[2117] & layer_0[7179]); 
    assign out[7811] = ~layer_0[186]; 
    assign out[7812] = ~(layer_0[7248] ^ layer_0[2495]); 
    assign out[7813] = layer_0[3696] & layer_0[1335]; 
    assign out[7814] = layer_0[415] ^ layer_0[10251]; 
    assign out[7815] = ~(layer_0[4028] | layer_0[3909]); 
    assign out[7816] = ~(layer_0[6050] ^ layer_0[6970]); 
    assign out[7817] = layer_0[7019]; 
    assign out[7818] = ~(layer_0[11380] ^ layer_0[6933]); 
    assign out[7819] = layer_0[11432] & ~layer_0[1832]; 
    assign out[7820] = ~layer_0[4992] | (layer_0[532] & layer_0[4992]); 
    assign out[7821] = layer_0[725] ^ layer_0[139]; 
    assign out[7822] = ~layer_0[11577]; 
    assign out[7823] = ~(layer_0[10805] ^ layer_0[1606]); 
    assign out[7824] = ~layer_0[7710]; 
    assign out[7825] = ~(layer_0[8892] ^ layer_0[9869]); 
    assign out[7826] = layer_0[11674]; 
    assign out[7827] = ~(layer_0[628] | layer_0[3624]); 
    assign out[7828] = layer_0[746] ^ layer_0[1727]; 
    assign out[7829] = layer_0[2366]; 
    assign out[7830] = layer_0[1984] ^ layer_0[9643]; 
    assign out[7831] = layer_0[3746] & ~layer_0[5442]; 
    assign out[7832] = ~(layer_0[9266] & layer_0[6109]); 
    assign out[7833] = layer_0[2747] ^ layer_0[5518]; 
    assign out[7834] = layer_0[7411] & layer_0[392]; 
    assign out[7835] = ~(layer_0[6027] ^ layer_0[1423]); 
    assign out[7836] = layer_0[6755] & layer_0[11453]; 
    assign out[7837] = layer_0[7437] & ~layer_0[8958]; 
    assign out[7838] = ~(layer_0[5956] ^ layer_0[11950]); 
    assign out[7839] = ~layer_0[82]; 
    assign out[7840] = layer_0[8161]; 
    assign out[7841] = layer_0[2314]; 
    assign out[7842] = layer_0[5650] & layer_0[9706]; 
    assign out[7843] = ~layer_0[5092] | (layer_0[5092] & layer_0[8025]); 
    assign out[7844] = ~(layer_0[919] ^ layer_0[5721]); 
    assign out[7845] = layer_0[718] & layer_0[5242]; 
    assign out[7846] = ~(layer_0[941] | layer_0[4359]); 
    assign out[7847] = ~layer_0[3381]; 
    assign out[7848] = layer_0[8358] | layer_0[4139]; 
    assign out[7849] = ~(layer_0[2295] ^ layer_0[137]); 
    assign out[7850] = ~(layer_0[11088] ^ layer_0[3118]); 
    assign out[7851] = ~(layer_0[11734] | layer_0[2046]); 
    assign out[7852] = ~layer_0[9857] | (layer_0[1127] & layer_0[9857]); 
    assign out[7853] = layer_0[8008] ^ layer_0[9854]; 
    assign out[7854] = layer_0[7911] & ~layer_0[1427]; 
    assign out[7855] = layer_0[7172] ^ layer_0[3800]; 
    assign out[7856] = ~(layer_0[6148] ^ layer_0[5440]); 
    assign out[7857] = layer_0[3672] ^ layer_0[2672]; 
    assign out[7858] = layer_0[4112] & layer_0[5290]; 
    assign out[7859] = ~(layer_0[4751] & layer_0[1295]); 
    assign out[7860] = ~layer_0[10826]; 
    assign out[7861] = ~(layer_0[3091] ^ layer_0[5993]); 
    assign out[7862] = layer_0[11603] & ~layer_0[2534]; 
    assign out[7863] = ~layer_0[4223]; 
    assign out[7864] = layer_0[11859] & ~layer_0[4842]; 
    assign out[7865] = ~(layer_0[11211] ^ layer_0[518]); 
    assign out[7866] = ~layer_0[8958]; 
    assign out[7867] = ~(layer_0[6333] | layer_0[3478]); 
    assign out[7868] = ~(layer_0[8460] ^ layer_0[5627]); 
    assign out[7869] = layer_0[8998] ^ layer_0[9866]; 
    assign out[7870] = ~(layer_0[10536] | layer_0[7273]); 
    assign out[7871] = ~(layer_0[5549] ^ layer_0[11678]); 
    assign out[7872] = layer_0[10764] ^ layer_0[4148]; 
    assign out[7873] = ~layer_0[2317]; 
    assign out[7874] = ~(layer_0[5228] ^ layer_0[9353]); 
    assign out[7875] = layer_0[9608]; 
    assign out[7876] = ~(layer_0[11347] ^ layer_0[2695]); 
    assign out[7877] = layer_0[3980] & ~layer_0[11673]; 
    assign out[7878] = ~(layer_0[5240] | layer_0[9511]); 
    assign out[7879] = layer_0[7887] ^ layer_0[10325]; 
    assign out[7880] = layer_0[3315]; 
    assign out[7881] = ~layer_0[1296]; 
    assign out[7882] = layer_0[10102]; 
    assign out[7883] = layer_0[11532] & ~layer_0[428]; 
    assign out[7884] = ~(layer_0[1578] | layer_0[5992]); 
    assign out[7885] = ~layer_0[3580]; 
    assign out[7886] = ~layer_0[8507]; 
    assign out[7887] = layer_0[7758] & ~layer_0[11331]; 
    assign out[7888] = layer_0[10265] & ~layer_0[6854]; 
    assign out[7889] = layer_0[6963] & layer_0[2927]; 
    assign out[7890] = layer_0[475] & layer_0[1826]; 
    assign out[7891] = layer_0[106] | layer_0[6731]; 
    assign out[7892] = layer_0[8251]; 
    assign out[7893] = layer_0[3295] & layer_0[11615]; 
    assign out[7894] = layer_0[6547] & ~layer_0[8899]; 
    assign out[7895] = ~(layer_0[352] | layer_0[5506]); 
    assign out[7896] = layer_0[1931] & layer_0[7540]; 
    assign out[7897] = layer_0[8026] & layer_0[11035]; 
    assign out[7898] = layer_0[7422]; 
    assign out[7899] = layer_0[1774]; 
    assign out[7900] = ~(layer_0[2772] | layer_0[7788]); 
    assign out[7901] = ~(layer_0[11681] | layer_0[10562]); 
    assign out[7902] = layer_0[4388] & layer_0[9795]; 
    assign out[7903] = ~(layer_0[9449] ^ layer_0[786]); 
    assign out[7904] = ~(layer_0[968] ^ layer_0[9429]); 
    assign out[7905] = ~layer_0[7063] | (layer_0[7063] & layer_0[1275]); 
    assign out[7906] = layer_0[8130] & ~layer_0[2546]; 
    assign out[7907] = layer_0[1842] | layer_0[4947]; 
    assign out[7908] = layer_0[7083] & ~layer_0[8933]; 
    assign out[7909] = ~(layer_0[2766] | layer_0[3608]); 
    assign out[7910] = layer_0[1381] & ~layer_0[750]; 
    assign out[7911] = layer_0[5761] & ~layer_0[11272]; 
    assign out[7912] = layer_0[11128] | layer_0[6031]; 
    assign out[7913] = ~(layer_0[11732] | layer_0[6472]); 
    assign out[7914] = ~(layer_0[11513] ^ layer_0[3722]); 
    assign out[7915] = ~(layer_0[918] ^ layer_0[9702]); 
    assign out[7916] = layer_0[4170] ^ layer_0[3123]; 
    assign out[7917] = layer_0[1253] & ~layer_0[9848]; 
    assign out[7918] = ~layer_0[10629] | (layer_0[10629] & layer_0[9950]); 
    assign out[7919] = ~(layer_0[11164] & layer_0[567]); 
    assign out[7920] = layer_0[4948] & ~layer_0[759]; 
    assign out[7921] = layer_0[2924]; 
    assign out[7922] = ~(layer_0[2638] | layer_0[11682]); 
    assign out[7923] = ~layer_0[267]; 
    assign out[7924] = layer_0[11688] ^ layer_0[2302]; 
    assign out[7925] = ~layer_0[7163]; 
    assign out[7926] = ~layer_0[6028]; 
    assign out[7927] = layer_0[11764] & layer_0[2315]; 
    assign out[7928] = ~layer_0[9169]; 
    assign out[7929] = layer_0[6409]; 
    assign out[7930] = layer_0[6769] ^ layer_0[7814]; 
    assign out[7931] = layer_0[9667]; 
    assign out[7932] = layer_0[7146] ^ layer_0[5118]; 
    assign out[7933] = ~layer_0[7988] | (layer_0[7988] & layer_0[10032]); 
    assign out[7934] = layer_0[8531] & ~layer_0[2537]; 
    assign out[7935] = ~(layer_0[5320] | layer_0[8800]); 
    assign out[7936] = layer_0[3207] & ~layer_0[123]; 
    assign out[7937] = ~(layer_0[4507] ^ layer_0[3321]); 
    assign out[7938] = layer_0[150] ^ layer_0[4077]; 
    assign out[7939] = ~(layer_0[4715] ^ layer_0[6556]); 
    assign out[7940] = ~(layer_0[602] | layer_0[8956]); 
    assign out[7941] = ~layer_0[630]; 
    assign out[7942] = layer_0[4248] & ~layer_0[9902]; 
    assign out[7943] = layer_0[2354] & layer_0[2535]; 
    assign out[7944] = layer_0[6820] & ~layer_0[4700]; 
    assign out[7945] = ~layer_0[961]; 
    assign out[7946] = ~(layer_0[121] & layer_0[1829]); 
    assign out[7947] = layer_0[9856] & layer_0[4771]; 
    assign out[7948] = layer_0[9593]; 
    assign out[7949] = layer_0[10310] & ~layer_0[2855]; 
    assign out[7950] = layer_0[94] ^ layer_0[6039]; 
    assign out[7951] = ~(layer_0[6655] ^ layer_0[10044]); 
    assign out[7952] = layer_0[7939]; 
    assign out[7953] = ~(layer_0[10666] | layer_0[6614]); 
    assign out[7954] = ~(layer_0[11136] ^ layer_0[11257]); 
    assign out[7955] = ~(layer_0[1286] & layer_0[4324]); 
    assign out[7956] = layer_0[8289] ^ layer_0[4059]; 
    assign out[7957] = ~layer_0[749]; 
    assign out[7958] = layer_0[4415] & ~layer_0[9315]; 
    assign out[7959] = ~(layer_0[1229] | layer_0[1757]); 
    assign out[7960] = layer_0[1946] & ~layer_0[8458]; 
    assign out[7961] = layer_0[596] & ~layer_0[2142]; 
    assign out[7962] = ~layer_0[10979] | (layer_0[10979] & layer_0[9013]); 
    assign out[7963] = ~layer_0[3705]; 
    assign out[7964] = layer_0[6843] & layer_0[6945]; 
    assign out[7965] = ~(layer_0[7759] | layer_0[6432]); 
    assign out[7966] = layer_0[1004] & layer_0[11582]; 
    assign out[7967] = layer_0[8254] | layer_0[6244]; 
    assign out[7968] = layer_0[8159] & layer_0[8531]; 
    assign out[7969] = ~(layer_0[4201] ^ layer_0[701]); 
    assign out[7970] = layer_0[10986]; 
    assign out[7971] = layer_0[3576]; 
    assign out[7972] = ~(layer_0[1496] ^ layer_0[10197]); 
    assign out[7973] = layer_0[4945] | layer_0[4398]; 
    assign out[7974] = ~(layer_0[5146] ^ layer_0[10616]); 
    assign out[7975] = layer_0[1250] ^ layer_0[7595]; 
    assign out[7976] = layer_0[4376]; 
    assign out[7977] = layer_0[4140] & ~layer_0[8817]; 
    assign out[7978] = ~(layer_0[325] | layer_0[11298]); 
    assign out[7979] = ~layer_0[6154]; 
    assign out[7980] = ~(layer_0[10294] & layer_0[5638]); 
    assign out[7981] = layer_0[838]; 
    assign out[7982] = layer_0[5210] & layer_0[10582]; 
    assign out[7983] = ~(layer_0[929] ^ layer_0[850]); 
    assign out[7984] = layer_0[9355] & ~layer_0[10506]; 
    assign out[7985] = ~layer_0[3143]; 
    assign out[7986] = ~(layer_0[4702] | layer_0[3390]); 
    assign out[7987] = ~(layer_0[1956] | layer_0[10523]); 
    assign out[7988] = layer_0[2792]; 
    assign out[7989] = ~(layer_0[11219] | layer_0[3681]); 
    assign out[7990] = layer_0[9824] ^ layer_0[3783]; 
    assign out[7991] = ~layer_0[18]; 
    assign out[7992] = layer_0[9396] & layer_0[1165]; 
    assign out[7993] = ~(layer_0[10360] ^ layer_0[2844]); 
    assign out[7994] = ~layer_0[6795] | (layer_0[6795] & layer_0[3151]); 
    assign out[7995] = layer_0[8903] & layer_0[4968]; 
    assign out[7996] = layer_0[2152] | layer_0[1291]; 
    assign out[7997] = layer_0[1463] & layer_0[1876]; 
    assign out[7998] = layer_0[2869] & ~layer_0[808]; 
    assign out[7999] = ~layer_0[4113]; 
    assign out[8000] = 1'b0; 
    assign out[8001] = 1'b0; 
    assign out[8002] = 1'b0; 
    assign out[8003] = 1'b0; 
    assign out[8004] = 1'b0; 
    assign out[8005] = 1'b0; 
    assign out[8006] = 1'b0; 
    assign out[8007] = 1'b0; 
    assign out[8008] = 1'b0; 
    assign out[8009] = 1'b0; 
    assign out[8010] = 1'b0; 
    assign out[8011] = 1'b0; 
    assign out[8012] = 1'b0; 
    assign out[8013] = 1'b0; 
    assign out[8014] = 1'b0; 
    assign out[8015] = 1'b0; 
    assign out[8016] = 1'b0; 
    assign out[8017] = 1'b0; 
    assign out[8018] = 1'b0; 
    assign out[8019] = 1'b0; 
    assign out[8020] = 1'b0; 
    assign out[8021] = 1'b0; 
    assign out[8022] = 1'b0; 
    assign out[8023] = 1'b0; 
    assign out[8024] = 1'b0; 
    assign out[8025] = 1'b0; 
    assign out[8026] = 1'b0; 
    assign out[8027] = 1'b0; 
    assign out[8028] = 1'b0; 
    assign out[8029] = 1'b0; 
    assign out[8030] = 1'b0; 
    assign out[8031] = 1'b0; 
    assign out[8032] = 1'b0; 
    assign out[8033] = 1'b0; 
    assign out[8034] = 1'b0; 
    assign out[8035] = 1'b0; 
    assign out[8036] = 1'b0; 
    assign out[8037] = 1'b0; 
    assign out[8038] = 1'b0; 
    assign out[8039] = 1'b0; 
    assign out[8040] = 1'b0; 
    assign out[8041] = 1'b0; 
    assign out[8042] = 1'b0; 
    assign out[8043] = 1'b0; 
    assign out[8044] = 1'b0; 
    assign out[8045] = 1'b0; 
    assign out[8046] = 1'b0; 
    assign out[8047] = 1'b0; 
    assign out[8048] = 1'b0; 
    assign out[8049] = 1'b0; 
    assign out[8050] = 1'b0; 
    assign out[8051] = 1'b0; 
    assign out[8052] = 1'b0; 
    assign out[8053] = 1'b0; 
    assign out[8054] = 1'b0; 
    assign out[8055] = 1'b0; 
    assign out[8056] = 1'b0; 
    assign out[8057] = 1'b0; 
    assign out[8058] = 1'b0; 
    assign out[8059] = 1'b0; 
    assign out[8060] = 1'b0; 
    assign out[8061] = 1'b0; 
    assign out[8062] = 1'b0; 
    assign out[8063] = 1'b0; 
    assign out[8064] = 1'b0; 
    assign out[8065] = 1'b0; 
    assign out[8066] = 1'b0; 
    assign out[8067] = 1'b0; 
    assign out[8068] = 1'b0; 
    assign out[8069] = 1'b0; 
    assign out[8070] = 1'b0; 
    assign out[8071] = 1'b0; 
    assign out[8072] = 1'b0; 
    assign out[8073] = 1'b0; 
    assign out[8074] = 1'b0; 
    assign out[8075] = 1'b0; 
    assign out[8076] = 1'b0; 
    assign out[8077] = 1'b0; 
    assign out[8078] = 1'b0; 
    assign out[8079] = 1'b0; 
    assign out[8080] = 1'b0; 
    assign out[8081] = 1'b0; 
    assign out[8082] = 1'b0; 
    assign out[8083] = 1'b0; 
    assign out[8084] = 1'b0; 
    assign out[8085] = 1'b0; 
    assign out[8086] = 1'b0; 
    assign out[8087] = 1'b0; 
    assign out[8088] = 1'b0; 
    assign out[8089] = 1'b0; 
    assign out[8090] = 1'b0; 
    assign out[8091] = 1'b0; 
    assign out[8092] = 1'b0; 
    assign out[8093] = 1'b0; 
    assign out[8094] = 1'b0; 
    assign out[8095] = 1'b0; 
    assign out[8096] = 1'b0; 
    assign out[8097] = 1'b0; 
    assign out[8098] = 1'b0; 
    assign out[8099] = 1'b0; 
    assign out[8100] = 1'b0; 
    assign out[8101] = 1'b0; 
    assign out[8102] = 1'b0; 
    assign out[8103] = 1'b0; 
    assign out[8104] = 1'b0; 
    assign out[8105] = 1'b0; 
    assign out[8106] = 1'b0; 
    assign out[8107] = 1'b0; 
    assign out[8108] = 1'b0; 
    assign out[8109] = 1'b0; 
    assign out[8110] = 1'b0; 
    assign out[8111] = 1'b0; 
    assign out[8112] = 1'b0; 
    assign out[8113] = 1'b0; 
    assign out[8114] = 1'b0; 
    assign out[8115] = 1'b0; 
    assign out[8116] = 1'b0; 
    assign out[8117] = 1'b0; 
    assign out[8118] = 1'b0; 
    assign out[8119] = 1'b0; 
    assign out[8120] = 1'b0; 
    assign out[8121] = 1'b0; 
    assign out[8122] = 1'b0; 
    assign out[8123] = 1'b0; 
    assign out[8124] = 1'b0; 
    assign out[8125] = 1'b0; 
    assign out[8126] = 1'b0; 
    assign out[8127] = 1'b0; 
    assign out[8128] = 1'b0; 
    assign out[8129] = 1'b0; 
    assign out[8130] = 1'b0; 
    assign out[8131] = 1'b0; 
    assign out[8132] = 1'b0; 
    assign out[8133] = 1'b0; 
    assign out[8134] = 1'b0; 
    assign out[8135] = 1'b0; 
    assign out[8136] = 1'b0; 
    assign out[8137] = 1'b0; 
    assign out[8138] = 1'b0; 
    assign out[8139] = 1'b0; 
    assign out[8140] = 1'b0; 
    assign out[8141] = 1'b0; 
    assign out[8142] = 1'b0; 
    assign out[8143] = 1'b0; 
    assign out[8144] = 1'b0; 
    assign out[8145] = 1'b0; 
    assign out[8146] = 1'b0; 
    assign out[8147] = 1'b0; 
    assign out[8148] = 1'b0; 
    assign out[8149] = 1'b0; 
    assign out[8150] = 1'b0; 
    assign out[8151] = 1'b0; 
    assign out[8152] = 1'b0; 
    assign out[8153] = 1'b0; 
    assign out[8154] = 1'b0; 
    assign out[8155] = 1'b0; 
    assign out[8156] = 1'b0; 
    assign out[8157] = 1'b0; 
    assign out[8158] = 1'b0; 
    assign out[8159] = 1'b0; 
    assign out[8160] = 1'b0; 
    assign out[8161] = 1'b0; 
    assign out[8162] = 1'b0; 
    assign out[8163] = 1'b0; 
    assign out[8164] = 1'b0; 
    assign out[8165] = 1'b0; 
    assign out[8166] = 1'b0; 
    assign out[8167] = 1'b0; 
    assign out[8168] = 1'b0; 
    assign out[8169] = 1'b0; 
    assign out[8170] = 1'b0; 
    assign out[8171] = 1'b0; 
    assign out[8172] = 1'b0; 
    assign out[8173] = 1'b0; 
    assign out[8174] = 1'b0; 
    assign out[8175] = 1'b0; 
    assign out[8176] = 1'b0; 
    assign out[8177] = 1'b0; 
    assign out[8178] = 1'b0; 
    assign out[8179] = 1'b0; 
    assign out[8180] = 1'b0; 
    assign out[8181] = 1'b0; 
    assign out[8182] = 1'b0; 
    assign out[8183] = 1'b0; 
    assign out[8184] = 1'b0; 
    assign out[8185] = 1'b0; 
    assign out[8186] = 1'b0; 
    assign out[8187] = 1'b0; 
    assign out[8188] = 1'b0; 
    assign out[8189] = 1'b0; 
    assign out[8190] = 1'b0; 
    assign out[8191] = 1'b0; 
    assign out[8192] = 1'b0; 
    assign out[8193] = 1'b0; 
    assign out[8194] = 1'b0; 
    assign out[8195] = 1'b0; 
    assign out[8196] = 1'b0; 
    assign out[8197] = 1'b0; 
    assign out[8198] = 1'b0; 
    assign out[8199] = 1'b0; 
    assign out[8200] = 1'b0; 
    assign out[8201] = 1'b0; 
    assign out[8202] = 1'b0; 
    assign out[8203] = 1'b0; 
    assign out[8204] = 1'b0; 
    assign out[8205] = 1'b0; 
    assign out[8206] = 1'b0; 
    assign out[8207] = 1'b0; 
    assign out[8208] = 1'b0; 
    assign out[8209] = 1'b0; 
    assign out[8210] = 1'b0; 
    assign out[8211] = 1'b0; 
    assign out[8212] = 1'b0; 
    assign out[8213] = 1'b0; 
    assign out[8214] = 1'b0; 
    assign out[8215] = 1'b0; 
    assign out[8216] = 1'b0; 
    assign out[8217] = 1'b0; 
    assign out[8218] = 1'b0; 
    assign out[8219] = 1'b0; 
    assign out[8220] = 1'b0; 
    assign out[8221] = 1'b0; 
    assign out[8222] = 1'b0; 
    assign out[8223] = 1'b0; 
    assign out[8224] = 1'b0; 
    assign out[8225] = 1'b0; 
    assign out[8226] = 1'b0; 
    assign out[8227] = 1'b0; 
    assign out[8228] = 1'b0; 
    assign out[8229] = 1'b0; 
    assign out[8230] = 1'b0; 
    assign out[8231] = 1'b0; 
    assign out[8232] = 1'b0; 
    assign out[8233] = 1'b0; 
    assign out[8234] = 1'b0; 
    assign out[8235] = 1'b0; 
    assign out[8236] = 1'b0; 
    assign out[8237] = 1'b0; 
    assign out[8238] = 1'b0; 
    assign out[8239] = 1'b0; 
    assign out[8240] = 1'b0; 
    assign out[8241] = 1'b0; 
    assign out[8242] = 1'b0; 
    assign out[8243] = 1'b0; 
    assign out[8244] = 1'b0; 
    assign out[8245] = 1'b0; 
    assign out[8246] = 1'b0; 
    assign out[8247] = 1'b0; 
    assign out[8248] = 1'b0; 
    assign out[8249] = 1'b0; 
    assign out[8250] = 1'b0; 
    assign out[8251] = 1'b0; 
    assign out[8252] = 1'b0; 
    assign out[8253] = 1'b0; 
    assign out[8254] = 1'b0; 
    assign out[8255] = 1'b0; 
    assign out[8256] = 1'b0; 
    assign out[8257] = 1'b0; 
    assign out[8258] = 1'b0; 
    assign out[8259] = 1'b0; 
    assign out[8260] = 1'b0; 
    assign out[8261] = 1'b0; 
    assign out[8262] = 1'b0; 
    assign out[8263] = 1'b0; 
    assign out[8264] = 1'b0; 
    assign out[8265] = 1'b0; 
    assign out[8266] = 1'b0; 
    assign out[8267] = 1'b0; 
    assign out[8268] = 1'b0; 
    assign out[8269] = 1'b0; 
    assign out[8270] = 1'b0; 
    assign out[8271] = 1'b0; 
    assign out[8272] = 1'b0; 
    assign out[8273] = 1'b0; 
    assign out[8274] = 1'b0; 
    assign out[8275] = 1'b0; 
    assign out[8276] = 1'b0; 
    assign out[8277] = 1'b0; 
    assign out[8278] = 1'b0; 
    assign out[8279] = 1'b0; 
    assign out[8280] = 1'b0; 
    assign out[8281] = 1'b0; 
    assign out[8282] = 1'b0; 
    assign out[8283] = 1'b0; 
    assign out[8284] = 1'b0; 
    assign out[8285] = 1'b0; 
    assign out[8286] = 1'b0; 
    assign out[8287] = 1'b0; 
    assign out[8288] = 1'b0; 
    assign out[8289] = 1'b0; 
    assign out[8290] = 1'b0; 
    assign out[8291] = 1'b0; 
    assign out[8292] = 1'b0; 
    assign out[8293] = 1'b0; 
    assign out[8294] = 1'b0; 
    assign out[8295] = 1'b0; 
    assign out[8296] = 1'b0; 
    assign out[8297] = 1'b0; 
    assign out[8298] = 1'b0; 
    assign out[8299] = 1'b0; 
    assign out[8300] = 1'b0; 
    assign out[8301] = 1'b0; 
    assign out[8302] = 1'b0; 
    assign out[8303] = 1'b0; 
    assign out[8304] = 1'b0; 
    assign out[8305] = 1'b0; 
    assign out[8306] = 1'b0; 
    assign out[8307] = 1'b0; 
    assign out[8308] = 1'b0; 
    assign out[8309] = 1'b0; 
    assign out[8310] = 1'b0; 
    assign out[8311] = 1'b0; 
    assign out[8312] = 1'b0; 
    assign out[8313] = 1'b0; 
    assign out[8314] = 1'b0; 
    assign out[8315] = 1'b0; 
    assign out[8316] = 1'b0; 
    assign out[8317] = 1'b0; 
    assign out[8318] = 1'b0; 
    assign out[8319] = 1'b0; 
    assign out[8320] = 1'b0; 
    assign out[8321] = 1'b0; 
    assign out[8322] = 1'b0; 
    assign out[8323] = 1'b0; 
    assign out[8324] = 1'b0; 
    assign out[8325] = 1'b0; 
    assign out[8326] = 1'b0; 
    assign out[8327] = 1'b0; 
    assign out[8328] = 1'b0; 
    assign out[8329] = 1'b0; 
    assign out[8330] = 1'b0; 
    assign out[8331] = 1'b0; 
    assign out[8332] = 1'b0; 
    assign out[8333] = 1'b0; 
    assign out[8334] = 1'b0; 
    assign out[8335] = 1'b0; 
    assign out[8336] = 1'b0; 
    assign out[8337] = 1'b0; 
    assign out[8338] = 1'b0; 
    assign out[8339] = 1'b0; 
    assign out[8340] = 1'b0; 
    assign out[8341] = 1'b0; 
    assign out[8342] = 1'b0; 
    assign out[8343] = 1'b0; 
    assign out[8344] = 1'b0; 
    assign out[8345] = 1'b0; 
    assign out[8346] = 1'b0; 
    assign out[8347] = 1'b0; 
    assign out[8348] = 1'b0; 
    assign out[8349] = 1'b0; 
    assign out[8350] = 1'b0; 
    assign out[8351] = 1'b0; 
    assign out[8352] = 1'b0; 
    assign out[8353] = 1'b0; 
    assign out[8354] = 1'b0; 
    assign out[8355] = 1'b0; 
    assign out[8356] = 1'b0; 
    assign out[8357] = 1'b0; 
    assign out[8358] = 1'b0; 
    assign out[8359] = 1'b0; 
    assign out[8360] = 1'b0; 
    assign out[8361] = 1'b0; 
    assign out[8362] = 1'b0; 
    assign out[8363] = 1'b0; 
    assign out[8364] = 1'b0; 
    assign out[8365] = 1'b0; 
    assign out[8366] = 1'b0; 
    assign out[8367] = 1'b0; 
    assign out[8368] = 1'b0; 
    assign out[8369] = 1'b0; 
    assign out[8370] = 1'b0; 
    assign out[8371] = 1'b0; 
    assign out[8372] = 1'b0; 
    assign out[8373] = 1'b0; 
    assign out[8374] = 1'b0; 
    assign out[8375] = 1'b0; 
    assign out[8376] = 1'b0; 
    assign out[8377] = 1'b0; 
    assign out[8378] = 1'b0; 
    assign out[8379] = 1'b0; 
    assign out[8380] = 1'b0; 
    assign out[8381] = 1'b0; 
    assign out[8382] = 1'b0; 
    assign out[8383] = 1'b0; 
    assign out[8384] = 1'b0; 
    assign out[8385] = 1'b0; 
    assign out[8386] = 1'b0; 
    assign out[8387] = 1'b0; 
    assign out[8388] = 1'b0; 
    assign out[8389] = 1'b0; 
    assign out[8390] = 1'b0; 
    assign out[8391] = 1'b0; 
    assign out[8392] = 1'b0; 
    assign out[8393] = 1'b0; 
    assign out[8394] = 1'b0; 
    assign out[8395] = 1'b0; 
    assign out[8396] = 1'b0; 
    assign out[8397] = 1'b0; 
    assign out[8398] = 1'b0; 
    assign out[8399] = 1'b0; 
    assign out[8400] = 1'b0; 
    assign out[8401] = 1'b0; 
    assign out[8402] = 1'b0; 
    assign out[8403] = 1'b0; 
    assign out[8404] = 1'b0; 
    assign out[8405] = 1'b0; 
    assign out[8406] = 1'b0; 
    assign out[8407] = 1'b0; 
    assign out[8408] = 1'b0; 
    assign out[8409] = 1'b0; 
    assign out[8410] = 1'b0; 
    assign out[8411] = 1'b0; 
    assign out[8412] = 1'b0; 
    assign out[8413] = 1'b0; 
    assign out[8414] = 1'b0; 
    assign out[8415] = 1'b0; 
    assign out[8416] = 1'b0; 
    assign out[8417] = 1'b0; 
    assign out[8418] = 1'b0; 
    assign out[8419] = 1'b0; 
    assign out[8420] = 1'b0; 
    assign out[8421] = 1'b0; 
    assign out[8422] = 1'b0; 
    assign out[8423] = 1'b0; 
    assign out[8424] = 1'b0; 
    assign out[8425] = 1'b0; 
    assign out[8426] = 1'b0; 
    assign out[8427] = 1'b0; 
    assign out[8428] = 1'b0; 
    assign out[8429] = 1'b0; 
    assign out[8430] = 1'b0; 
    assign out[8431] = 1'b0; 
    assign out[8432] = 1'b0; 
    assign out[8433] = 1'b0; 
    assign out[8434] = 1'b0; 
    assign out[8435] = 1'b0; 
    assign out[8436] = 1'b0; 
    assign out[8437] = 1'b0; 
    assign out[8438] = 1'b0; 
    assign out[8439] = 1'b0; 
    assign out[8440] = 1'b0; 
    assign out[8441] = 1'b0; 
    assign out[8442] = 1'b0; 
    assign out[8443] = 1'b0; 
    assign out[8444] = 1'b0; 
    assign out[8445] = 1'b0; 
    assign out[8446] = 1'b0; 
    assign out[8447] = 1'b0; 
    assign out[8448] = 1'b0; 
    assign out[8449] = 1'b0; 
    assign out[8450] = 1'b0; 
    assign out[8451] = 1'b0; 
    assign out[8452] = 1'b0; 
    assign out[8453] = 1'b0; 
    assign out[8454] = 1'b0; 
    assign out[8455] = 1'b0; 
    assign out[8456] = 1'b0; 
    assign out[8457] = 1'b0; 
    assign out[8458] = 1'b0; 
    assign out[8459] = 1'b0; 
    assign out[8460] = 1'b0; 
    assign out[8461] = 1'b0; 
    assign out[8462] = 1'b0; 
    assign out[8463] = 1'b0; 
    assign out[8464] = 1'b0; 
    assign out[8465] = 1'b0; 
    assign out[8466] = 1'b0; 
    assign out[8467] = 1'b0; 
    assign out[8468] = 1'b0; 
    assign out[8469] = 1'b0; 
    assign out[8470] = 1'b0; 
    assign out[8471] = 1'b0; 
    assign out[8472] = 1'b0; 
    assign out[8473] = 1'b0; 
    assign out[8474] = 1'b0; 
    assign out[8475] = 1'b0; 
    assign out[8476] = 1'b0; 
    assign out[8477] = 1'b0; 
    assign out[8478] = 1'b0; 
    assign out[8479] = 1'b0; 
    assign out[8480] = 1'b0; 
    assign out[8481] = 1'b0; 
    assign out[8482] = 1'b0; 
    assign out[8483] = 1'b0; 
    assign out[8484] = 1'b0; 
    assign out[8485] = 1'b0; 
    assign out[8486] = 1'b0; 
    assign out[8487] = 1'b0; 
    assign out[8488] = 1'b0; 
    assign out[8489] = 1'b0; 
    assign out[8490] = 1'b0; 
    assign out[8491] = 1'b0; 
    assign out[8492] = 1'b0; 
    assign out[8493] = 1'b0; 
    assign out[8494] = 1'b0; 
    assign out[8495] = 1'b0; 
    assign out[8496] = 1'b0; 
    assign out[8497] = 1'b0; 
    assign out[8498] = 1'b0; 
    assign out[8499] = 1'b0; 
    assign out[8500] = 1'b0; 
    assign out[8501] = 1'b0; 
    assign out[8502] = 1'b0; 
    assign out[8503] = 1'b0; 
    assign out[8504] = 1'b0; 
    assign out[8505] = 1'b0; 
    assign out[8506] = 1'b0; 
    assign out[8507] = 1'b0; 
    assign out[8508] = 1'b0; 
    assign out[8509] = 1'b0; 
    assign out[8510] = 1'b0; 
    assign out[8511] = 1'b0; 
    assign out[8512] = 1'b0; 
    assign out[8513] = 1'b0; 
    assign out[8514] = 1'b0; 
    assign out[8515] = 1'b0; 
    assign out[8516] = 1'b0; 
    assign out[8517] = 1'b0; 
    assign out[8518] = 1'b0; 
    assign out[8519] = 1'b0; 
    assign out[8520] = 1'b0; 
    assign out[8521] = 1'b0; 
    assign out[8522] = 1'b0; 
    assign out[8523] = 1'b0; 
    assign out[8524] = 1'b0; 
    assign out[8525] = 1'b0; 
    assign out[8526] = 1'b0; 
    assign out[8527] = 1'b0; 
    assign out[8528] = 1'b0; 
    assign out[8529] = 1'b0; 
    assign out[8530] = 1'b0; 
    assign out[8531] = 1'b0; 
    assign out[8532] = 1'b0; 
    assign out[8533] = 1'b0; 
    assign out[8534] = 1'b0; 
    assign out[8535] = 1'b0; 
    assign out[8536] = 1'b0; 
    assign out[8537] = 1'b0; 
    assign out[8538] = 1'b0; 
    assign out[8539] = 1'b0; 
    assign out[8540] = 1'b0; 
    assign out[8541] = 1'b0; 
    assign out[8542] = 1'b0; 
    assign out[8543] = 1'b0; 
    assign out[8544] = 1'b0; 
    assign out[8545] = 1'b0; 
    assign out[8546] = 1'b0; 
    assign out[8547] = 1'b0; 
    assign out[8548] = 1'b0; 
    assign out[8549] = 1'b0; 
    assign out[8550] = 1'b0; 
    assign out[8551] = 1'b0; 
    assign out[8552] = 1'b0; 
    assign out[8553] = 1'b0; 
    assign out[8554] = 1'b0; 
    assign out[8555] = 1'b0; 
    assign out[8556] = 1'b0; 
    assign out[8557] = 1'b0; 
    assign out[8558] = 1'b0; 
    assign out[8559] = 1'b0; 
    assign out[8560] = 1'b0; 
    assign out[8561] = 1'b0; 
    assign out[8562] = 1'b0; 
    assign out[8563] = 1'b0; 
    assign out[8564] = 1'b0; 
    assign out[8565] = 1'b0; 
    assign out[8566] = 1'b0; 
    assign out[8567] = 1'b0; 
    assign out[8568] = 1'b0; 
    assign out[8569] = 1'b0; 
    assign out[8570] = 1'b0; 
    assign out[8571] = 1'b0; 
    assign out[8572] = 1'b0; 
    assign out[8573] = 1'b0; 
    assign out[8574] = 1'b0; 
    assign out[8575] = 1'b0; 
    assign out[8576] = 1'b0; 
    assign out[8577] = 1'b0; 
    assign out[8578] = 1'b0; 
    assign out[8579] = 1'b0; 
    assign out[8580] = 1'b0; 
    assign out[8581] = 1'b0; 
    assign out[8582] = 1'b0; 
    assign out[8583] = 1'b0; 
    assign out[8584] = 1'b0; 
    assign out[8585] = 1'b0; 
    assign out[8586] = 1'b0; 
    assign out[8587] = 1'b0; 
    assign out[8588] = 1'b0; 
    assign out[8589] = 1'b0; 
    assign out[8590] = 1'b0; 
    assign out[8591] = 1'b0; 
    assign out[8592] = 1'b0; 
    assign out[8593] = 1'b0; 
    assign out[8594] = 1'b0; 
    assign out[8595] = 1'b0; 
    assign out[8596] = 1'b0; 
    assign out[8597] = 1'b0; 
    assign out[8598] = 1'b0; 
    assign out[8599] = 1'b0; 
    assign out[8600] = 1'b0; 
    assign out[8601] = 1'b0; 
    assign out[8602] = 1'b0; 
    assign out[8603] = 1'b0; 
    assign out[8604] = 1'b0; 
    assign out[8605] = 1'b0; 
    assign out[8606] = 1'b0; 
    assign out[8607] = 1'b0; 
    assign out[8608] = 1'b0; 
    assign out[8609] = 1'b0; 
    assign out[8610] = 1'b0; 
    assign out[8611] = 1'b0; 
    assign out[8612] = 1'b0; 
    assign out[8613] = 1'b0; 
    assign out[8614] = 1'b0; 
    assign out[8615] = 1'b0; 
    assign out[8616] = 1'b0; 
    assign out[8617] = 1'b0; 
    assign out[8618] = 1'b0; 
    assign out[8619] = 1'b0; 
    assign out[8620] = 1'b0; 
    assign out[8621] = 1'b0; 
    assign out[8622] = 1'b0; 
    assign out[8623] = 1'b0; 
    assign out[8624] = 1'b0; 
    assign out[8625] = 1'b0; 
    assign out[8626] = 1'b0; 
    assign out[8627] = 1'b0; 
    assign out[8628] = 1'b0; 
    assign out[8629] = 1'b0; 
    assign out[8630] = 1'b0; 
    assign out[8631] = 1'b0; 
    assign out[8632] = 1'b0; 
    assign out[8633] = 1'b0; 
    assign out[8634] = 1'b0; 
    assign out[8635] = 1'b0; 
    assign out[8636] = 1'b0; 
    assign out[8637] = 1'b0; 
    assign out[8638] = 1'b0; 
    assign out[8639] = 1'b0; 
    assign out[8640] = 1'b0; 
    assign out[8641] = 1'b0; 
    assign out[8642] = 1'b0; 
    assign out[8643] = 1'b0; 
    assign out[8644] = 1'b0; 
    assign out[8645] = 1'b0; 
    assign out[8646] = 1'b0; 
    assign out[8647] = 1'b0; 
    assign out[8648] = 1'b0; 
    assign out[8649] = 1'b0; 
    assign out[8650] = 1'b0; 
    assign out[8651] = 1'b0; 
    assign out[8652] = 1'b0; 
    assign out[8653] = 1'b0; 
    assign out[8654] = 1'b0; 
    assign out[8655] = 1'b0; 
    assign out[8656] = 1'b0; 
    assign out[8657] = 1'b0; 
    assign out[8658] = 1'b0; 
    assign out[8659] = 1'b0; 
    assign out[8660] = 1'b0; 
    assign out[8661] = 1'b0; 
    assign out[8662] = 1'b0; 
    assign out[8663] = 1'b0; 
    assign out[8664] = 1'b0; 
    assign out[8665] = 1'b0; 
    assign out[8666] = 1'b0; 
    assign out[8667] = 1'b0; 
    assign out[8668] = 1'b0; 
    assign out[8669] = 1'b0; 
    assign out[8670] = 1'b0; 
    assign out[8671] = 1'b0; 
    assign out[8672] = 1'b0; 
    assign out[8673] = 1'b0; 
    assign out[8674] = 1'b0; 
    assign out[8675] = 1'b0; 
    assign out[8676] = 1'b0; 
    assign out[8677] = 1'b0; 
    assign out[8678] = 1'b0; 
    assign out[8679] = 1'b0; 
    assign out[8680] = 1'b0; 
    assign out[8681] = 1'b0; 
    assign out[8682] = 1'b0; 
    assign out[8683] = 1'b0; 
    assign out[8684] = 1'b0; 
    assign out[8685] = 1'b0; 
    assign out[8686] = 1'b0; 
    assign out[8687] = 1'b0; 
    assign out[8688] = 1'b0; 
    assign out[8689] = 1'b0; 
    assign out[8690] = 1'b0; 
    assign out[8691] = 1'b0; 
    assign out[8692] = 1'b0; 
    assign out[8693] = 1'b0; 
    assign out[8694] = 1'b0; 
    assign out[8695] = 1'b0; 
    assign out[8696] = 1'b0; 
    assign out[8697] = 1'b0; 
    assign out[8698] = 1'b0; 
    assign out[8699] = 1'b0; 
    assign out[8700] = 1'b0; 
    assign out[8701] = 1'b0; 
    assign out[8702] = 1'b0; 
    assign out[8703] = 1'b0; 
    assign out[8704] = 1'b0; 
    assign out[8705] = 1'b0; 
    assign out[8706] = 1'b0; 
    assign out[8707] = 1'b0; 
    assign out[8708] = 1'b0; 
    assign out[8709] = 1'b0; 
    assign out[8710] = 1'b0; 
    assign out[8711] = 1'b0; 
    assign out[8712] = 1'b0; 
    assign out[8713] = 1'b0; 
    assign out[8714] = 1'b0; 
    assign out[8715] = 1'b0; 
    assign out[8716] = 1'b0; 
    assign out[8717] = 1'b0; 
    assign out[8718] = 1'b0; 
    assign out[8719] = 1'b0; 
    assign out[8720] = 1'b0; 
    assign out[8721] = 1'b0; 
    assign out[8722] = 1'b0; 
    assign out[8723] = 1'b0; 
    assign out[8724] = 1'b0; 
    assign out[8725] = 1'b0; 
    assign out[8726] = 1'b0; 
    assign out[8727] = 1'b0; 
    assign out[8728] = 1'b0; 
    assign out[8729] = 1'b0; 
    assign out[8730] = 1'b0; 
    assign out[8731] = 1'b0; 
    assign out[8732] = 1'b0; 
    assign out[8733] = 1'b0; 
    assign out[8734] = 1'b0; 
    assign out[8735] = 1'b0; 
    assign out[8736] = 1'b0; 
    assign out[8737] = 1'b0; 
    assign out[8738] = 1'b0; 
    assign out[8739] = 1'b0; 
    assign out[8740] = 1'b0; 
    assign out[8741] = 1'b0; 
    assign out[8742] = 1'b0; 
    assign out[8743] = 1'b0; 
    assign out[8744] = 1'b0; 
    assign out[8745] = 1'b0; 
    assign out[8746] = 1'b0; 
    assign out[8747] = 1'b0; 
    assign out[8748] = 1'b0; 
    assign out[8749] = 1'b0; 
    assign out[8750] = 1'b0; 
    assign out[8751] = 1'b0; 
    assign out[8752] = 1'b0; 
    assign out[8753] = 1'b0; 
    assign out[8754] = 1'b0; 
    assign out[8755] = 1'b0; 
    assign out[8756] = 1'b0; 
    assign out[8757] = 1'b0; 
    assign out[8758] = 1'b0; 
    assign out[8759] = 1'b0; 
    assign out[8760] = 1'b0; 
    assign out[8761] = 1'b0; 
    assign out[8762] = 1'b0; 
    assign out[8763] = 1'b0; 
    assign out[8764] = 1'b0; 
    assign out[8765] = 1'b0; 
    assign out[8766] = 1'b0; 
    assign out[8767] = 1'b0; 
    assign out[8768] = 1'b0; 
    assign out[8769] = 1'b0; 
    assign out[8770] = 1'b0; 
    assign out[8771] = 1'b0; 
    assign out[8772] = 1'b0; 
    assign out[8773] = 1'b0; 
    assign out[8774] = 1'b0; 
    assign out[8775] = 1'b0; 
    assign out[8776] = 1'b0; 
    assign out[8777] = 1'b0; 
    assign out[8778] = 1'b0; 
    assign out[8779] = 1'b0; 
    assign out[8780] = 1'b0; 
    assign out[8781] = 1'b0; 
    assign out[8782] = 1'b0; 
    assign out[8783] = 1'b0; 
    assign out[8784] = 1'b0; 
    assign out[8785] = 1'b0; 
    assign out[8786] = 1'b0; 
    assign out[8787] = 1'b0; 
    assign out[8788] = 1'b0; 
    assign out[8789] = 1'b0; 
    assign out[8790] = 1'b0; 
    assign out[8791] = 1'b0; 
    assign out[8792] = 1'b0; 
    assign out[8793] = 1'b0; 
    assign out[8794] = 1'b0; 
    assign out[8795] = 1'b0; 
    assign out[8796] = 1'b0; 
    assign out[8797] = 1'b0; 
    assign out[8798] = 1'b0; 
    assign out[8799] = 1'b0; 
    assign out[8800] = 1'b0; 
    assign out[8801] = 1'b0; 
    assign out[8802] = 1'b0; 
    assign out[8803] = 1'b0; 
    assign out[8804] = 1'b0; 
    assign out[8805] = 1'b0; 
    assign out[8806] = 1'b0; 
    assign out[8807] = 1'b0; 
    assign out[8808] = 1'b0; 
    assign out[8809] = 1'b0; 
    assign out[8810] = 1'b0; 
    assign out[8811] = 1'b0; 
    assign out[8812] = 1'b0; 
    assign out[8813] = 1'b0; 
    assign out[8814] = 1'b0; 
    assign out[8815] = 1'b0; 
    assign out[8816] = 1'b0; 
    assign out[8817] = 1'b0; 
    assign out[8818] = 1'b0; 
    assign out[8819] = 1'b0; 
    assign out[8820] = 1'b0; 
    assign out[8821] = 1'b0; 
    assign out[8822] = 1'b0; 
    assign out[8823] = 1'b0; 
    assign out[8824] = 1'b0; 
    assign out[8825] = 1'b0; 
    assign out[8826] = 1'b0; 
    assign out[8827] = 1'b0; 
    assign out[8828] = 1'b0; 
    assign out[8829] = 1'b0; 
    assign out[8830] = 1'b0; 
    assign out[8831] = 1'b0; 
    assign out[8832] = 1'b0; 
    assign out[8833] = 1'b0; 
    assign out[8834] = 1'b0; 
    assign out[8835] = 1'b0; 
    assign out[8836] = 1'b0; 
    assign out[8837] = 1'b0; 
    assign out[8838] = 1'b0; 
    assign out[8839] = 1'b0; 
    assign out[8840] = 1'b0; 
    assign out[8841] = 1'b0; 
    assign out[8842] = 1'b0; 
    assign out[8843] = 1'b0; 
    assign out[8844] = 1'b0; 
    assign out[8845] = 1'b0; 
    assign out[8846] = 1'b0; 
    assign out[8847] = 1'b0; 
    assign out[8848] = 1'b0; 
    assign out[8849] = 1'b0; 
    assign out[8850] = 1'b0; 
    assign out[8851] = 1'b0; 
    assign out[8852] = 1'b0; 
    assign out[8853] = 1'b0; 
    assign out[8854] = 1'b0; 
    assign out[8855] = 1'b0; 
    assign out[8856] = 1'b0; 
    assign out[8857] = 1'b0; 
    assign out[8858] = 1'b0; 
    assign out[8859] = 1'b0; 
    assign out[8860] = 1'b0; 
    assign out[8861] = 1'b0; 
    assign out[8862] = 1'b0; 
    assign out[8863] = 1'b0; 
    assign out[8864] = 1'b0; 
    assign out[8865] = 1'b0; 
    assign out[8866] = 1'b0; 
    assign out[8867] = 1'b0; 
    assign out[8868] = 1'b0; 
    assign out[8869] = 1'b0; 
    assign out[8870] = 1'b0; 
    assign out[8871] = 1'b0; 
    assign out[8872] = 1'b0; 
    assign out[8873] = 1'b0; 
    assign out[8874] = 1'b0; 
    assign out[8875] = 1'b0; 
    assign out[8876] = 1'b0; 
    assign out[8877] = 1'b0; 
    assign out[8878] = 1'b0; 
    assign out[8879] = 1'b0; 
    assign out[8880] = 1'b0; 
    assign out[8881] = 1'b0; 
    assign out[8882] = 1'b0; 
    assign out[8883] = 1'b0; 
    assign out[8884] = 1'b0; 
    assign out[8885] = 1'b0; 
    assign out[8886] = 1'b0; 
    assign out[8887] = 1'b0; 
    assign out[8888] = 1'b0; 
    assign out[8889] = 1'b0; 
    assign out[8890] = 1'b0; 
    assign out[8891] = 1'b0; 
    assign out[8892] = 1'b0; 
    assign out[8893] = 1'b0; 
    assign out[8894] = 1'b0; 
    assign out[8895] = 1'b0; 
    assign out[8896] = 1'b0; 
    assign out[8897] = 1'b0; 
    assign out[8898] = 1'b0; 
    assign out[8899] = 1'b0; 
    assign out[8900] = 1'b0; 
    assign out[8901] = 1'b0; 
    assign out[8902] = 1'b0; 
    assign out[8903] = 1'b0; 
    assign out[8904] = 1'b0; 
    assign out[8905] = 1'b0; 
    assign out[8906] = 1'b0; 
    assign out[8907] = 1'b0; 
    assign out[8908] = 1'b0; 
    assign out[8909] = 1'b0; 
    assign out[8910] = 1'b0; 
    assign out[8911] = 1'b0; 
    assign out[8912] = 1'b0; 
    assign out[8913] = 1'b0; 
    assign out[8914] = 1'b0; 
    assign out[8915] = 1'b0; 
    assign out[8916] = 1'b0; 
    assign out[8917] = 1'b0; 
    assign out[8918] = 1'b0; 
    assign out[8919] = 1'b0; 
    assign out[8920] = 1'b0; 
    assign out[8921] = 1'b0; 
    assign out[8922] = 1'b0; 
    assign out[8923] = 1'b0; 
    assign out[8924] = 1'b0; 
    assign out[8925] = 1'b0; 
    assign out[8926] = 1'b0; 
    assign out[8927] = 1'b0; 
    assign out[8928] = 1'b0; 
    assign out[8929] = 1'b0; 
    assign out[8930] = 1'b0; 
    assign out[8931] = 1'b0; 
    assign out[8932] = 1'b0; 
    assign out[8933] = 1'b0; 
    assign out[8934] = 1'b0; 
    assign out[8935] = 1'b0; 
    assign out[8936] = 1'b0; 
    assign out[8937] = 1'b0; 
    assign out[8938] = 1'b0; 
    assign out[8939] = 1'b0; 
    assign out[8940] = 1'b0; 
    assign out[8941] = 1'b0; 
    assign out[8942] = 1'b0; 
    assign out[8943] = 1'b0; 
    assign out[8944] = 1'b0; 
    assign out[8945] = 1'b0; 
    assign out[8946] = 1'b0; 
    assign out[8947] = 1'b0; 
    assign out[8948] = 1'b0; 
    assign out[8949] = 1'b0; 
    assign out[8950] = 1'b0; 
    assign out[8951] = 1'b0; 
    assign out[8952] = 1'b0; 
    assign out[8953] = 1'b0; 
    assign out[8954] = 1'b0; 
    assign out[8955] = 1'b0; 
    assign out[8956] = 1'b0; 
    assign out[8957] = 1'b0; 
    assign out[8958] = 1'b0; 
    assign out[8959] = 1'b0; 
    assign out[8960] = 1'b0; 
    assign out[8961] = 1'b0; 
    assign out[8962] = 1'b0; 
    assign out[8963] = 1'b0; 
    assign out[8964] = 1'b0; 
    assign out[8965] = 1'b0; 
    assign out[8966] = 1'b0; 
    assign out[8967] = 1'b0; 
    assign out[8968] = 1'b0; 
    assign out[8969] = 1'b0; 
    assign out[8970] = 1'b0; 
    assign out[8971] = 1'b0; 
    assign out[8972] = 1'b0; 
    assign out[8973] = 1'b0; 
    assign out[8974] = 1'b0; 
    assign out[8975] = 1'b0; 
    assign out[8976] = 1'b0; 
    assign out[8977] = 1'b0; 
    assign out[8978] = 1'b0; 
    assign out[8979] = 1'b0; 
    assign out[8980] = 1'b0; 
    assign out[8981] = 1'b0; 
    assign out[8982] = 1'b0; 
    assign out[8983] = 1'b0; 
    assign out[8984] = 1'b0; 
    assign out[8985] = 1'b0; 
    assign out[8986] = 1'b0; 
    assign out[8987] = 1'b0; 
    assign out[8988] = 1'b0; 
    assign out[8989] = 1'b0; 
    assign out[8990] = 1'b0; 
    assign out[8991] = 1'b0; 
    assign out[8992] = 1'b0; 
    assign out[8993] = 1'b0; 
    assign out[8994] = 1'b0; 
    assign out[8995] = 1'b0; 
    assign out[8996] = 1'b0; 
    assign out[8997] = 1'b0; 
    assign out[8998] = 1'b0; 
    assign out[8999] = 1'b0; 
    assign out[9000] = 1'b0; 
    assign out[9001] = 1'b0; 
    assign out[9002] = 1'b0; 
    assign out[9003] = 1'b0; 
    assign out[9004] = 1'b0; 
    assign out[9005] = 1'b0; 
    assign out[9006] = 1'b0; 
    assign out[9007] = 1'b0; 
    assign out[9008] = 1'b0; 
    assign out[9009] = 1'b0; 
    assign out[9010] = 1'b0; 
    assign out[9011] = 1'b0; 
    assign out[9012] = 1'b0; 
    assign out[9013] = 1'b0; 
    assign out[9014] = 1'b0; 
    assign out[9015] = 1'b0; 
    assign out[9016] = 1'b0; 
    assign out[9017] = 1'b0; 
    assign out[9018] = 1'b0; 
    assign out[9019] = 1'b0; 
    assign out[9020] = 1'b0; 
    assign out[9021] = 1'b0; 
    assign out[9022] = 1'b0; 
    assign out[9023] = 1'b0; 
    assign out[9024] = 1'b0; 
    assign out[9025] = 1'b0; 
    assign out[9026] = 1'b0; 
    assign out[9027] = 1'b0; 
    assign out[9028] = 1'b0; 
    assign out[9029] = 1'b0; 
    assign out[9030] = 1'b0; 
    assign out[9031] = 1'b0; 
    assign out[9032] = 1'b0; 
    assign out[9033] = 1'b0; 
    assign out[9034] = 1'b0; 
    assign out[9035] = 1'b0; 
    assign out[9036] = 1'b0; 
    assign out[9037] = 1'b0; 
    assign out[9038] = 1'b0; 
    assign out[9039] = 1'b0; 
    assign out[9040] = 1'b0; 
    assign out[9041] = 1'b0; 
    assign out[9042] = 1'b0; 
    assign out[9043] = 1'b0; 
    assign out[9044] = 1'b0; 
    assign out[9045] = 1'b0; 
    assign out[9046] = 1'b0; 
    assign out[9047] = 1'b0; 
    assign out[9048] = 1'b0; 
    assign out[9049] = 1'b0; 
    assign out[9050] = 1'b0; 
    assign out[9051] = 1'b0; 
    assign out[9052] = 1'b0; 
    assign out[9053] = 1'b0; 
    assign out[9054] = 1'b0; 
    assign out[9055] = 1'b0; 
    assign out[9056] = 1'b0; 
    assign out[9057] = 1'b0; 
    assign out[9058] = 1'b0; 
    assign out[9059] = 1'b0; 
    assign out[9060] = 1'b0; 
    assign out[9061] = 1'b0; 
    assign out[9062] = 1'b0; 
    assign out[9063] = 1'b0; 
    assign out[9064] = 1'b0; 
    assign out[9065] = 1'b0; 
    assign out[9066] = 1'b0; 
    assign out[9067] = 1'b0; 
    assign out[9068] = 1'b0; 
    assign out[9069] = 1'b0; 
    assign out[9070] = 1'b0; 
    assign out[9071] = 1'b0; 
    assign out[9072] = 1'b0; 
    assign out[9073] = 1'b0; 
    assign out[9074] = 1'b0; 
    assign out[9075] = 1'b0; 
    assign out[9076] = 1'b0; 
    assign out[9077] = 1'b0; 
    assign out[9078] = 1'b0; 
    assign out[9079] = 1'b0; 
    assign out[9080] = 1'b0; 
    assign out[9081] = 1'b0; 
    assign out[9082] = 1'b0; 
    assign out[9083] = 1'b0; 
    assign out[9084] = 1'b0; 
    assign out[9085] = 1'b0; 
    assign out[9086] = 1'b0; 
    assign out[9087] = 1'b0; 
    assign out[9088] = 1'b0; 
    assign out[9089] = 1'b0; 
    assign out[9090] = 1'b0; 
    assign out[9091] = 1'b0; 
    assign out[9092] = 1'b0; 
    assign out[9093] = 1'b0; 
    assign out[9094] = 1'b0; 
    assign out[9095] = 1'b0; 
    assign out[9096] = 1'b0; 
    assign out[9097] = 1'b0; 
    assign out[9098] = 1'b0; 
    assign out[9099] = 1'b0; 
    assign out[9100] = 1'b0; 
    assign out[9101] = 1'b0; 
    assign out[9102] = 1'b0; 
    assign out[9103] = 1'b0; 
    assign out[9104] = 1'b0; 
    assign out[9105] = 1'b0; 
    assign out[9106] = 1'b0; 
    assign out[9107] = 1'b0; 
    assign out[9108] = 1'b0; 
    assign out[9109] = 1'b0; 
    assign out[9110] = 1'b0; 
    assign out[9111] = 1'b0; 
    assign out[9112] = 1'b0; 
    assign out[9113] = 1'b0; 
    assign out[9114] = 1'b0; 
    assign out[9115] = 1'b0; 
    assign out[9116] = 1'b0; 
    assign out[9117] = 1'b0; 
    assign out[9118] = 1'b0; 
    assign out[9119] = 1'b0; 
    assign out[9120] = 1'b0; 
    assign out[9121] = 1'b0; 
    assign out[9122] = 1'b0; 
    assign out[9123] = 1'b0; 
    assign out[9124] = 1'b0; 
    assign out[9125] = 1'b0; 
    assign out[9126] = 1'b0; 
    assign out[9127] = 1'b0; 
    assign out[9128] = 1'b0; 
    assign out[9129] = 1'b0; 
    assign out[9130] = 1'b0; 
    assign out[9131] = 1'b0; 
    assign out[9132] = 1'b0; 
    assign out[9133] = 1'b0; 
    assign out[9134] = 1'b0; 
    assign out[9135] = 1'b0; 
    assign out[9136] = 1'b0; 
    assign out[9137] = 1'b0; 
    assign out[9138] = 1'b0; 
    assign out[9139] = 1'b0; 
    assign out[9140] = 1'b0; 
    assign out[9141] = 1'b0; 
    assign out[9142] = 1'b0; 
    assign out[9143] = 1'b0; 
    assign out[9144] = 1'b0; 
    assign out[9145] = 1'b0; 
    assign out[9146] = 1'b0; 
    assign out[9147] = 1'b0; 
    assign out[9148] = 1'b0; 
    assign out[9149] = 1'b0; 
    assign out[9150] = 1'b0; 
    assign out[9151] = 1'b0; 
    assign out[9152] = 1'b0; 
    assign out[9153] = 1'b0; 
    assign out[9154] = 1'b0; 
    assign out[9155] = 1'b0; 
    assign out[9156] = 1'b0; 
    assign out[9157] = 1'b0; 
    assign out[9158] = 1'b0; 
    assign out[9159] = 1'b0; 
    assign out[9160] = 1'b0; 
    assign out[9161] = 1'b0; 
    assign out[9162] = 1'b0; 
    assign out[9163] = 1'b0; 
    assign out[9164] = 1'b0; 
    assign out[9165] = 1'b0; 
    assign out[9166] = 1'b0; 
    assign out[9167] = 1'b0; 
    assign out[9168] = 1'b0; 
    assign out[9169] = 1'b0; 
    assign out[9170] = 1'b0; 
    assign out[9171] = 1'b0; 
    assign out[9172] = 1'b0; 
    assign out[9173] = 1'b0; 
    assign out[9174] = 1'b0; 
    assign out[9175] = 1'b0; 
    assign out[9176] = 1'b0; 
    assign out[9177] = 1'b0; 
    assign out[9178] = 1'b0; 
    assign out[9179] = 1'b0; 
    assign out[9180] = 1'b0; 
    assign out[9181] = 1'b0; 
    assign out[9182] = 1'b0; 
    assign out[9183] = 1'b0; 
    assign out[9184] = 1'b0; 
    assign out[9185] = 1'b0; 
    assign out[9186] = 1'b0; 
    assign out[9187] = 1'b0; 
    assign out[9188] = 1'b0; 
    assign out[9189] = 1'b0; 
    assign out[9190] = 1'b0; 
    assign out[9191] = 1'b0; 
    assign out[9192] = 1'b0; 
    assign out[9193] = 1'b0; 
    assign out[9194] = 1'b0; 
    assign out[9195] = 1'b0; 
    assign out[9196] = 1'b0; 
    assign out[9197] = 1'b0; 
    assign out[9198] = 1'b0; 
    assign out[9199] = 1'b0; 
    assign out[9200] = 1'b0; 
    assign out[9201] = 1'b0; 
    assign out[9202] = 1'b0; 
    assign out[9203] = 1'b0; 
    assign out[9204] = 1'b0; 
    assign out[9205] = 1'b0; 
    assign out[9206] = 1'b0; 
    assign out[9207] = 1'b0; 
    assign out[9208] = 1'b0; 
    assign out[9209] = 1'b0; 
    assign out[9210] = 1'b0; 
    assign out[9211] = 1'b0; 
    assign out[9212] = 1'b0; 
    assign out[9213] = 1'b0; 
    assign out[9214] = 1'b0; 
    assign out[9215] = 1'b0; 
    assign out[9216] = 1'b0; 
    assign out[9217] = 1'b0; 
    assign out[9218] = 1'b0; 
    assign out[9219] = 1'b0; 
    assign out[9220] = 1'b0; 
    assign out[9221] = 1'b0; 
    assign out[9222] = 1'b0; 
    assign out[9223] = 1'b0; 
    assign out[9224] = 1'b0; 
    assign out[9225] = 1'b0; 
    assign out[9226] = 1'b0; 
    assign out[9227] = 1'b0; 
    assign out[9228] = 1'b0; 
    assign out[9229] = 1'b0; 
    assign out[9230] = 1'b0; 
    assign out[9231] = 1'b0; 
    assign out[9232] = 1'b0; 
    assign out[9233] = 1'b0; 
    assign out[9234] = 1'b0; 
    assign out[9235] = 1'b0; 
    assign out[9236] = 1'b0; 
    assign out[9237] = 1'b0; 
    assign out[9238] = 1'b0; 
    assign out[9239] = 1'b0; 
    assign out[9240] = 1'b0; 
    assign out[9241] = 1'b0; 
    assign out[9242] = 1'b0; 
    assign out[9243] = 1'b0; 
    assign out[9244] = 1'b0; 
    assign out[9245] = 1'b0; 
    assign out[9246] = 1'b0; 
    assign out[9247] = 1'b0; 
    assign out[9248] = 1'b0; 
    assign out[9249] = 1'b0; 
    assign out[9250] = 1'b0; 
    assign out[9251] = 1'b0; 
    assign out[9252] = 1'b0; 
    assign out[9253] = 1'b0; 
    assign out[9254] = 1'b0; 
    assign out[9255] = 1'b0; 
    assign out[9256] = 1'b0; 
    assign out[9257] = 1'b0; 
    assign out[9258] = 1'b0; 
    assign out[9259] = 1'b0; 
    assign out[9260] = 1'b0; 
    assign out[9261] = 1'b0; 
    assign out[9262] = 1'b0; 
    assign out[9263] = 1'b0; 
    assign out[9264] = 1'b0; 
    assign out[9265] = 1'b0; 
    assign out[9266] = 1'b0; 
    assign out[9267] = 1'b0; 
    assign out[9268] = 1'b0; 
    assign out[9269] = 1'b0; 
    assign out[9270] = 1'b0; 
    assign out[9271] = 1'b0; 
    assign out[9272] = 1'b0; 
    assign out[9273] = 1'b0; 
    assign out[9274] = 1'b0; 
    assign out[9275] = 1'b0; 
    assign out[9276] = 1'b0; 
    assign out[9277] = 1'b0; 
    assign out[9278] = 1'b0; 
    assign out[9279] = 1'b0; 
    assign out[9280] = 1'b0; 
    assign out[9281] = 1'b0; 
    assign out[9282] = 1'b0; 
    assign out[9283] = 1'b0; 
    assign out[9284] = 1'b0; 
    assign out[9285] = 1'b0; 
    assign out[9286] = 1'b0; 
    assign out[9287] = 1'b0; 
    assign out[9288] = 1'b0; 
    assign out[9289] = 1'b0; 
    assign out[9290] = 1'b0; 
    assign out[9291] = 1'b0; 
    assign out[9292] = 1'b0; 
    assign out[9293] = 1'b0; 
    assign out[9294] = 1'b0; 
    assign out[9295] = 1'b0; 
    assign out[9296] = 1'b0; 
    assign out[9297] = 1'b0; 
    assign out[9298] = 1'b0; 
    assign out[9299] = 1'b0; 
    assign out[9300] = 1'b0; 
    assign out[9301] = 1'b0; 
    assign out[9302] = 1'b0; 
    assign out[9303] = 1'b0; 
    assign out[9304] = 1'b0; 
    assign out[9305] = 1'b0; 
    assign out[9306] = 1'b0; 
    assign out[9307] = 1'b0; 
    assign out[9308] = 1'b0; 
    assign out[9309] = 1'b0; 
    assign out[9310] = 1'b0; 
    assign out[9311] = 1'b0; 
    assign out[9312] = 1'b0; 
    assign out[9313] = 1'b0; 
    assign out[9314] = 1'b0; 
    assign out[9315] = 1'b0; 
    assign out[9316] = 1'b0; 
    assign out[9317] = 1'b0; 
    assign out[9318] = 1'b0; 
    assign out[9319] = 1'b0; 
    assign out[9320] = 1'b0; 
    assign out[9321] = 1'b0; 
    assign out[9322] = 1'b0; 
    assign out[9323] = 1'b0; 
    assign out[9324] = 1'b0; 
    assign out[9325] = 1'b0; 
    assign out[9326] = 1'b0; 
    assign out[9327] = 1'b0; 
    assign out[9328] = 1'b0; 
    assign out[9329] = 1'b0; 
    assign out[9330] = 1'b0; 
    assign out[9331] = 1'b0; 
    assign out[9332] = 1'b0; 
    assign out[9333] = 1'b0; 
    assign out[9334] = 1'b0; 
    assign out[9335] = 1'b0; 
    assign out[9336] = 1'b0; 
    assign out[9337] = 1'b0; 
    assign out[9338] = 1'b0; 
    assign out[9339] = 1'b0; 
    assign out[9340] = 1'b0; 
    assign out[9341] = 1'b0; 
    assign out[9342] = 1'b0; 
    assign out[9343] = 1'b0; 
    assign out[9344] = 1'b0; 
    assign out[9345] = 1'b0; 
    assign out[9346] = 1'b0; 
    assign out[9347] = 1'b0; 
    assign out[9348] = 1'b0; 
    assign out[9349] = 1'b0; 
    assign out[9350] = 1'b0; 
    assign out[9351] = 1'b0; 
    assign out[9352] = 1'b0; 
    assign out[9353] = 1'b0; 
    assign out[9354] = 1'b0; 
    assign out[9355] = 1'b0; 
    assign out[9356] = 1'b0; 
    assign out[9357] = 1'b0; 
    assign out[9358] = 1'b0; 
    assign out[9359] = 1'b0; 
    assign out[9360] = 1'b0; 
    assign out[9361] = 1'b0; 
    assign out[9362] = 1'b0; 
    assign out[9363] = 1'b0; 
    assign out[9364] = 1'b0; 
    assign out[9365] = 1'b0; 
    assign out[9366] = 1'b0; 
    assign out[9367] = 1'b0; 
    assign out[9368] = 1'b0; 
    assign out[9369] = 1'b0; 
    assign out[9370] = 1'b0; 
    assign out[9371] = 1'b0; 
    assign out[9372] = 1'b0; 
    assign out[9373] = 1'b0; 
    assign out[9374] = 1'b0; 
    assign out[9375] = 1'b0; 
    assign out[9376] = 1'b0; 
    assign out[9377] = 1'b0; 
    assign out[9378] = 1'b0; 
    assign out[9379] = 1'b0; 
    assign out[9380] = 1'b0; 
    assign out[9381] = 1'b0; 
    assign out[9382] = 1'b0; 
    assign out[9383] = 1'b0; 
    assign out[9384] = 1'b0; 
    assign out[9385] = 1'b0; 
    assign out[9386] = 1'b0; 
    assign out[9387] = 1'b0; 
    assign out[9388] = 1'b0; 
    assign out[9389] = 1'b0; 
    assign out[9390] = 1'b0; 
    assign out[9391] = 1'b0; 
    assign out[9392] = 1'b0; 
    assign out[9393] = 1'b0; 
    assign out[9394] = 1'b0; 
    assign out[9395] = 1'b0; 
    assign out[9396] = 1'b0; 
    assign out[9397] = 1'b0; 
    assign out[9398] = 1'b0; 
    assign out[9399] = 1'b0; 
    assign out[9400] = 1'b0; 
    assign out[9401] = 1'b0; 
    assign out[9402] = 1'b0; 
    assign out[9403] = 1'b0; 
    assign out[9404] = 1'b0; 
    assign out[9405] = 1'b0; 
    assign out[9406] = 1'b0; 
    assign out[9407] = 1'b0; 
    assign out[9408] = 1'b0; 
    assign out[9409] = 1'b0; 
    assign out[9410] = 1'b0; 
    assign out[9411] = 1'b0; 
    assign out[9412] = 1'b0; 
    assign out[9413] = 1'b0; 
    assign out[9414] = 1'b0; 
    assign out[9415] = 1'b0; 
    assign out[9416] = 1'b0; 
    assign out[9417] = 1'b0; 
    assign out[9418] = 1'b0; 
    assign out[9419] = 1'b0; 
    assign out[9420] = 1'b0; 
    assign out[9421] = 1'b0; 
    assign out[9422] = 1'b0; 
    assign out[9423] = 1'b0; 
    assign out[9424] = 1'b0; 
    assign out[9425] = 1'b0; 
    assign out[9426] = 1'b0; 
    assign out[9427] = 1'b0; 
    assign out[9428] = 1'b0; 
    assign out[9429] = 1'b0; 
    assign out[9430] = 1'b0; 
    assign out[9431] = 1'b0; 
    assign out[9432] = 1'b0; 
    assign out[9433] = 1'b0; 
    assign out[9434] = 1'b0; 
    assign out[9435] = 1'b0; 
    assign out[9436] = 1'b0; 
    assign out[9437] = 1'b0; 
    assign out[9438] = 1'b0; 
    assign out[9439] = 1'b0; 
    assign out[9440] = 1'b0; 
    assign out[9441] = 1'b0; 
    assign out[9442] = 1'b0; 
    assign out[9443] = 1'b0; 
    assign out[9444] = 1'b0; 
    assign out[9445] = 1'b0; 
    assign out[9446] = 1'b0; 
    assign out[9447] = 1'b0; 
    assign out[9448] = 1'b0; 
    assign out[9449] = 1'b0; 
    assign out[9450] = 1'b0; 
    assign out[9451] = 1'b0; 
    assign out[9452] = 1'b0; 
    assign out[9453] = 1'b0; 
    assign out[9454] = 1'b0; 
    assign out[9455] = 1'b0; 
    assign out[9456] = 1'b0; 
    assign out[9457] = 1'b0; 
    assign out[9458] = 1'b0; 
    assign out[9459] = 1'b0; 
    assign out[9460] = 1'b0; 
    assign out[9461] = 1'b0; 
    assign out[9462] = 1'b0; 
    assign out[9463] = 1'b0; 
    assign out[9464] = 1'b0; 
    assign out[9465] = 1'b0; 
    assign out[9466] = 1'b0; 
    assign out[9467] = 1'b0; 
    assign out[9468] = 1'b0; 
    assign out[9469] = 1'b0; 
    assign out[9470] = 1'b0; 
    assign out[9471] = 1'b0; 
    assign out[9472] = 1'b0; 
    assign out[9473] = 1'b0; 
    assign out[9474] = 1'b0; 
    assign out[9475] = 1'b0; 
    assign out[9476] = 1'b0; 
    assign out[9477] = 1'b0; 
    assign out[9478] = 1'b0; 
    assign out[9479] = 1'b0; 
    assign out[9480] = 1'b0; 
    assign out[9481] = 1'b0; 
    assign out[9482] = 1'b0; 
    assign out[9483] = 1'b0; 
    assign out[9484] = 1'b0; 
    assign out[9485] = 1'b0; 
    assign out[9486] = 1'b0; 
    assign out[9487] = 1'b0; 
    assign out[9488] = 1'b0; 
    assign out[9489] = 1'b0; 
    assign out[9490] = 1'b0; 
    assign out[9491] = 1'b0; 
    assign out[9492] = 1'b0; 
    assign out[9493] = 1'b0; 
    assign out[9494] = 1'b0; 
    assign out[9495] = 1'b0; 
    assign out[9496] = 1'b0; 
    assign out[9497] = 1'b0; 
    assign out[9498] = 1'b0; 
    assign out[9499] = 1'b0; 
    assign out[9500] = 1'b0; 
    assign out[9501] = 1'b0; 
    assign out[9502] = 1'b0; 
    assign out[9503] = 1'b0; 
    assign out[9504] = 1'b0; 
    assign out[9505] = 1'b0; 
    assign out[9506] = 1'b0; 
    assign out[9507] = 1'b0; 
    assign out[9508] = 1'b0; 
    assign out[9509] = 1'b0; 
    assign out[9510] = 1'b0; 
    assign out[9511] = 1'b0; 
    assign out[9512] = 1'b0; 
    assign out[9513] = 1'b0; 
    assign out[9514] = 1'b0; 
    assign out[9515] = 1'b0; 
    assign out[9516] = 1'b0; 
    assign out[9517] = 1'b0; 
    assign out[9518] = 1'b0; 
    assign out[9519] = 1'b0; 
    assign out[9520] = 1'b0; 
    assign out[9521] = 1'b0; 
    assign out[9522] = 1'b0; 
    assign out[9523] = 1'b0; 
    assign out[9524] = 1'b0; 
    assign out[9525] = 1'b0; 
    assign out[9526] = 1'b0; 
    assign out[9527] = 1'b0; 
    assign out[9528] = 1'b0; 
    assign out[9529] = 1'b0; 
    assign out[9530] = 1'b0; 
    assign out[9531] = 1'b0; 
    assign out[9532] = 1'b0; 
    assign out[9533] = 1'b0; 
    assign out[9534] = 1'b0; 
    assign out[9535] = 1'b0; 
    assign out[9536] = 1'b0; 
    assign out[9537] = 1'b0; 
    assign out[9538] = 1'b0; 
    assign out[9539] = 1'b0; 
    assign out[9540] = 1'b0; 
    assign out[9541] = 1'b0; 
    assign out[9542] = 1'b0; 
    assign out[9543] = 1'b0; 
    assign out[9544] = 1'b0; 
    assign out[9545] = 1'b0; 
    assign out[9546] = 1'b0; 
    assign out[9547] = 1'b0; 
    assign out[9548] = 1'b0; 
    assign out[9549] = 1'b0; 
    assign out[9550] = 1'b0; 
    assign out[9551] = 1'b0; 
    assign out[9552] = 1'b0; 
    assign out[9553] = 1'b0; 
    assign out[9554] = 1'b0; 
    assign out[9555] = 1'b0; 
    assign out[9556] = 1'b0; 
    assign out[9557] = 1'b0; 
    assign out[9558] = 1'b0; 
    assign out[9559] = 1'b0; 
    assign out[9560] = 1'b0; 
    assign out[9561] = 1'b0; 
    assign out[9562] = 1'b0; 
    assign out[9563] = 1'b0; 
    assign out[9564] = 1'b0; 
    assign out[9565] = 1'b0; 
    assign out[9566] = 1'b0; 
    assign out[9567] = 1'b0; 
    assign out[9568] = 1'b0; 
    assign out[9569] = 1'b0; 
    assign out[9570] = 1'b0; 
    assign out[9571] = 1'b0; 
    assign out[9572] = 1'b0; 
    assign out[9573] = 1'b0; 
    assign out[9574] = 1'b0; 
    assign out[9575] = 1'b0; 
    assign out[9576] = 1'b0; 
    assign out[9577] = 1'b0; 
    assign out[9578] = 1'b0; 
    assign out[9579] = 1'b0; 
    assign out[9580] = 1'b0; 
    assign out[9581] = 1'b0; 
    assign out[9582] = 1'b0; 
    assign out[9583] = 1'b0; 
    assign out[9584] = 1'b0; 
    assign out[9585] = 1'b0; 
    assign out[9586] = 1'b0; 
    assign out[9587] = 1'b0; 
    assign out[9588] = 1'b0; 
    assign out[9589] = 1'b0; 
    assign out[9590] = 1'b0; 
    assign out[9591] = 1'b0; 
    assign out[9592] = 1'b0; 
    assign out[9593] = 1'b0; 
    assign out[9594] = 1'b0; 
    assign out[9595] = 1'b0; 
    assign out[9596] = 1'b0; 
    assign out[9597] = 1'b0; 
    assign out[9598] = 1'b0; 
    assign out[9599] = 1'b0; 
    assign out[9600] = 1'b0; 
    assign out[9601] = 1'b0; 
    assign out[9602] = 1'b0; 
    assign out[9603] = 1'b0; 
    assign out[9604] = 1'b0; 
    assign out[9605] = 1'b0; 
    assign out[9606] = 1'b0; 
    assign out[9607] = 1'b0; 
    assign out[9608] = 1'b0; 
    assign out[9609] = 1'b0; 
    assign out[9610] = 1'b0; 
    assign out[9611] = 1'b0; 
    assign out[9612] = 1'b0; 
    assign out[9613] = 1'b0; 
    assign out[9614] = 1'b0; 
    assign out[9615] = 1'b0; 
    assign out[9616] = 1'b0; 
    assign out[9617] = 1'b0; 
    assign out[9618] = 1'b0; 
    assign out[9619] = 1'b0; 
    assign out[9620] = 1'b0; 
    assign out[9621] = 1'b0; 
    assign out[9622] = 1'b0; 
    assign out[9623] = 1'b0; 
    assign out[9624] = 1'b0; 
    assign out[9625] = 1'b0; 
    assign out[9626] = 1'b0; 
    assign out[9627] = 1'b0; 
    assign out[9628] = 1'b0; 
    assign out[9629] = 1'b0; 
    assign out[9630] = 1'b0; 
    assign out[9631] = 1'b0; 
    assign out[9632] = 1'b0; 
    assign out[9633] = 1'b0; 
    assign out[9634] = 1'b0; 
    assign out[9635] = 1'b0; 
    assign out[9636] = 1'b0; 
    assign out[9637] = 1'b0; 
    assign out[9638] = 1'b0; 
    assign out[9639] = 1'b0; 
    assign out[9640] = 1'b0; 
    assign out[9641] = 1'b0; 
    assign out[9642] = 1'b0; 
    assign out[9643] = 1'b0; 
    assign out[9644] = 1'b0; 
    assign out[9645] = 1'b0; 
    assign out[9646] = 1'b0; 
    assign out[9647] = 1'b0; 
    assign out[9648] = 1'b0; 
    assign out[9649] = 1'b0; 
    assign out[9650] = 1'b0; 
    assign out[9651] = 1'b0; 
    assign out[9652] = 1'b0; 
    assign out[9653] = 1'b0; 
    assign out[9654] = 1'b0; 
    assign out[9655] = 1'b0; 
    assign out[9656] = 1'b0; 
    assign out[9657] = 1'b0; 
    assign out[9658] = 1'b0; 
    assign out[9659] = 1'b0; 
    assign out[9660] = 1'b0; 
    assign out[9661] = 1'b0; 
    assign out[9662] = 1'b0; 
    assign out[9663] = 1'b0; 
    assign out[9664] = 1'b0; 
    assign out[9665] = 1'b0; 
    assign out[9666] = 1'b0; 
    assign out[9667] = 1'b0; 
    assign out[9668] = 1'b0; 
    assign out[9669] = 1'b0; 
    assign out[9670] = 1'b0; 
    assign out[9671] = 1'b0; 
    assign out[9672] = 1'b0; 
    assign out[9673] = 1'b0; 
    assign out[9674] = 1'b0; 
    assign out[9675] = 1'b0; 
    assign out[9676] = 1'b0; 
    assign out[9677] = 1'b0; 
    assign out[9678] = 1'b0; 
    assign out[9679] = 1'b0; 
    assign out[9680] = 1'b0; 
    assign out[9681] = 1'b0; 
    assign out[9682] = 1'b0; 
    assign out[9683] = 1'b0; 
    assign out[9684] = 1'b0; 
    assign out[9685] = 1'b0; 
    assign out[9686] = 1'b0; 
    assign out[9687] = 1'b0; 
    assign out[9688] = 1'b0; 
    assign out[9689] = 1'b0; 
    assign out[9690] = 1'b0; 
    assign out[9691] = 1'b0; 
    assign out[9692] = 1'b0; 
    assign out[9693] = 1'b0; 
    assign out[9694] = 1'b0; 
    assign out[9695] = 1'b0; 
    assign out[9696] = 1'b0; 
    assign out[9697] = 1'b0; 
    assign out[9698] = 1'b0; 
    assign out[9699] = 1'b0; 
    assign out[9700] = 1'b0; 
    assign out[9701] = 1'b0; 
    assign out[9702] = 1'b0; 
    assign out[9703] = 1'b0; 
    assign out[9704] = 1'b0; 
    assign out[9705] = 1'b0; 
    assign out[9706] = 1'b0; 
    assign out[9707] = 1'b0; 
    assign out[9708] = 1'b0; 
    assign out[9709] = 1'b0; 
    assign out[9710] = 1'b0; 
    assign out[9711] = 1'b0; 
    assign out[9712] = 1'b0; 
    assign out[9713] = 1'b0; 
    assign out[9714] = 1'b0; 
    assign out[9715] = 1'b0; 
    assign out[9716] = 1'b0; 
    assign out[9717] = 1'b0; 
    assign out[9718] = 1'b0; 
    assign out[9719] = 1'b0; 
    assign out[9720] = 1'b0; 
    assign out[9721] = 1'b0; 
    assign out[9722] = 1'b0; 
    assign out[9723] = 1'b0; 
    assign out[9724] = 1'b0; 
    assign out[9725] = 1'b0; 
    assign out[9726] = 1'b0; 
    assign out[9727] = 1'b0; 
    assign out[9728] = 1'b0; 
    assign out[9729] = 1'b0; 
    assign out[9730] = 1'b0; 
    assign out[9731] = 1'b0; 
    assign out[9732] = 1'b0; 
    assign out[9733] = 1'b0; 
    assign out[9734] = 1'b0; 
    assign out[9735] = 1'b0; 
    assign out[9736] = 1'b0; 
    assign out[9737] = 1'b0; 
    assign out[9738] = 1'b0; 
    assign out[9739] = 1'b0; 
    assign out[9740] = 1'b0; 
    assign out[9741] = 1'b0; 
    assign out[9742] = 1'b0; 
    assign out[9743] = 1'b0; 
    assign out[9744] = 1'b0; 
    assign out[9745] = 1'b0; 
    assign out[9746] = 1'b0; 
    assign out[9747] = 1'b0; 
    assign out[9748] = 1'b0; 
    assign out[9749] = 1'b0; 
    assign out[9750] = 1'b0; 
    assign out[9751] = 1'b0; 
    assign out[9752] = 1'b0; 
    assign out[9753] = 1'b0; 
    assign out[9754] = 1'b0; 
    assign out[9755] = 1'b0; 
    assign out[9756] = 1'b0; 
    assign out[9757] = 1'b0; 
    assign out[9758] = 1'b0; 
    assign out[9759] = 1'b0; 
    assign out[9760] = 1'b0; 
    assign out[9761] = 1'b0; 
    assign out[9762] = 1'b0; 
    assign out[9763] = 1'b0; 
    assign out[9764] = 1'b0; 
    assign out[9765] = 1'b0; 
    assign out[9766] = 1'b0; 
    assign out[9767] = 1'b0; 
    assign out[9768] = 1'b0; 
    assign out[9769] = 1'b0; 
    assign out[9770] = 1'b0; 
    assign out[9771] = 1'b0; 
    assign out[9772] = 1'b0; 
    assign out[9773] = 1'b0; 
    assign out[9774] = 1'b0; 
    assign out[9775] = 1'b0; 
    assign out[9776] = 1'b0; 
    assign out[9777] = 1'b0; 
    assign out[9778] = 1'b0; 
    assign out[9779] = 1'b0; 
    assign out[9780] = 1'b0; 
    assign out[9781] = 1'b0; 
    assign out[9782] = 1'b0; 
    assign out[9783] = 1'b0; 
    assign out[9784] = 1'b0; 
    assign out[9785] = 1'b0; 
    assign out[9786] = 1'b0; 
    assign out[9787] = 1'b0; 
    assign out[9788] = 1'b0; 
    assign out[9789] = 1'b0; 
    assign out[9790] = 1'b0; 
    assign out[9791] = 1'b0; 
    assign out[9792] = 1'b0; 
    assign out[9793] = 1'b0; 
    assign out[9794] = 1'b0; 
    assign out[9795] = 1'b0; 
    assign out[9796] = 1'b0; 
    assign out[9797] = 1'b0; 
    assign out[9798] = 1'b0; 
    assign out[9799] = 1'b0; 
    assign out[9800] = 1'b0; 
    assign out[9801] = 1'b0; 
    assign out[9802] = 1'b0; 
    assign out[9803] = 1'b0; 
    assign out[9804] = 1'b0; 
    assign out[9805] = 1'b0; 
    assign out[9806] = 1'b0; 
    assign out[9807] = 1'b0; 
    assign out[9808] = 1'b0; 
    assign out[9809] = 1'b0; 
    assign out[9810] = 1'b0; 
    assign out[9811] = 1'b0; 
    assign out[9812] = 1'b0; 
    assign out[9813] = 1'b0; 
    assign out[9814] = 1'b0; 
    assign out[9815] = 1'b0; 
    assign out[9816] = 1'b0; 
    assign out[9817] = 1'b0; 
    assign out[9818] = 1'b0; 
    assign out[9819] = 1'b0; 
    assign out[9820] = 1'b0; 
    assign out[9821] = 1'b0; 
    assign out[9822] = 1'b0; 
    assign out[9823] = 1'b0; 
    assign out[9824] = 1'b0; 
    assign out[9825] = 1'b0; 
    assign out[9826] = 1'b0; 
    assign out[9827] = 1'b0; 
    assign out[9828] = 1'b0; 
    assign out[9829] = 1'b0; 
    assign out[9830] = 1'b0; 
    assign out[9831] = 1'b0; 
    assign out[9832] = 1'b0; 
    assign out[9833] = 1'b0; 
    assign out[9834] = 1'b0; 
    assign out[9835] = 1'b0; 
    assign out[9836] = 1'b0; 
    assign out[9837] = 1'b0; 
    assign out[9838] = 1'b0; 
    assign out[9839] = 1'b0; 
    assign out[9840] = 1'b0; 
    assign out[9841] = 1'b0; 
    assign out[9842] = 1'b0; 
    assign out[9843] = 1'b0; 
    assign out[9844] = 1'b0; 
    assign out[9845] = 1'b0; 
    assign out[9846] = 1'b0; 
    assign out[9847] = 1'b0; 
    assign out[9848] = 1'b0; 
    assign out[9849] = 1'b0; 
    assign out[9850] = 1'b0; 
    assign out[9851] = 1'b0; 
    assign out[9852] = 1'b0; 
    assign out[9853] = 1'b0; 
    assign out[9854] = 1'b0; 
    assign out[9855] = 1'b0; 
    assign out[9856] = 1'b0; 
    assign out[9857] = 1'b0; 
    assign out[9858] = 1'b0; 
    assign out[9859] = 1'b0; 
    assign out[9860] = 1'b0; 
    assign out[9861] = 1'b0; 
    assign out[9862] = 1'b0; 
    assign out[9863] = 1'b0; 
    assign out[9864] = 1'b0; 
    assign out[9865] = 1'b0; 
    assign out[9866] = 1'b0; 
    assign out[9867] = 1'b0; 
    assign out[9868] = 1'b0; 
    assign out[9869] = 1'b0; 
    assign out[9870] = 1'b0; 
    assign out[9871] = 1'b0; 
    assign out[9872] = 1'b0; 
    assign out[9873] = 1'b0; 
    assign out[9874] = 1'b0; 
    assign out[9875] = 1'b0; 
    assign out[9876] = 1'b0; 
    assign out[9877] = 1'b0; 
    assign out[9878] = 1'b0; 
    assign out[9879] = 1'b0; 
    assign out[9880] = 1'b0; 
    assign out[9881] = 1'b0; 
    assign out[9882] = 1'b0; 
    assign out[9883] = 1'b0; 
    assign out[9884] = 1'b0; 
    assign out[9885] = 1'b0; 
    assign out[9886] = 1'b0; 
    assign out[9887] = 1'b0; 
    assign out[9888] = 1'b0; 
    assign out[9889] = 1'b0; 
    assign out[9890] = 1'b0; 
    assign out[9891] = 1'b0; 
    assign out[9892] = 1'b0; 
    assign out[9893] = 1'b0; 
    assign out[9894] = 1'b0; 
    assign out[9895] = 1'b0; 
    assign out[9896] = 1'b0; 
    assign out[9897] = 1'b0; 
    assign out[9898] = 1'b0; 
    assign out[9899] = 1'b0; 
    assign out[9900] = 1'b0; 
    assign out[9901] = 1'b0; 
    assign out[9902] = 1'b0; 
    assign out[9903] = 1'b0; 
    assign out[9904] = 1'b0; 
    assign out[9905] = 1'b0; 
    assign out[9906] = 1'b0; 
    assign out[9907] = 1'b0; 
    assign out[9908] = 1'b0; 
    assign out[9909] = 1'b0; 
    assign out[9910] = 1'b0; 
    assign out[9911] = 1'b0; 
    assign out[9912] = 1'b0; 
    assign out[9913] = 1'b0; 
    assign out[9914] = 1'b0; 
    assign out[9915] = 1'b0; 
    assign out[9916] = 1'b0; 
    assign out[9917] = 1'b0; 
    assign out[9918] = 1'b0; 
    assign out[9919] = 1'b0; 
    assign out[9920] = 1'b0; 
    assign out[9921] = 1'b0; 
    assign out[9922] = 1'b0; 
    assign out[9923] = 1'b0; 
    assign out[9924] = 1'b0; 
    assign out[9925] = 1'b0; 
    assign out[9926] = 1'b0; 
    assign out[9927] = 1'b0; 
    assign out[9928] = 1'b0; 
    assign out[9929] = 1'b0; 
    assign out[9930] = 1'b0; 
    assign out[9931] = 1'b0; 
    assign out[9932] = 1'b0; 
    assign out[9933] = 1'b0; 
    assign out[9934] = 1'b0; 
    assign out[9935] = 1'b0; 
    assign out[9936] = 1'b0; 
    assign out[9937] = 1'b0; 
    assign out[9938] = 1'b0; 
    assign out[9939] = 1'b0; 
    assign out[9940] = 1'b0; 
    assign out[9941] = 1'b0; 
    assign out[9942] = 1'b0; 
    assign out[9943] = 1'b0; 
    assign out[9944] = 1'b0; 
    assign out[9945] = 1'b0; 
    assign out[9946] = 1'b0; 
    assign out[9947] = 1'b0; 
    assign out[9948] = 1'b0; 
    assign out[9949] = 1'b0; 
    assign out[9950] = 1'b0; 
    assign out[9951] = 1'b0; 
    assign out[9952] = 1'b0; 
    assign out[9953] = 1'b0; 
    assign out[9954] = 1'b0; 
    assign out[9955] = 1'b0; 
    assign out[9956] = 1'b0; 
    assign out[9957] = 1'b0; 
    assign out[9958] = 1'b0; 
    assign out[9959] = 1'b0; 
    assign out[9960] = 1'b0; 
    assign out[9961] = 1'b0; 
    assign out[9962] = 1'b0; 
    assign out[9963] = 1'b0; 
    assign out[9964] = 1'b0; 
    assign out[9965] = 1'b0; 
    assign out[9966] = 1'b0; 
    assign out[9967] = 1'b0; 
    assign out[9968] = 1'b0; 
    assign out[9969] = 1'b0; 
    assign out[9970] = 1'b0; 
    assign out[9971] = 1'b0; 
    assign out[9972] = 1'b0; 
    assign out[9973] = 1'b0; 
    assign out[9974] = 1'b0; 
    assign out[9975] = 1'b0; 
    assign out[9976] = 1'b0; 
    assign out[9977] = 1'b0; 
    assign out[9978] = 1'b0; 
    assign out[9979] = 1'b0; 
    assign out[9980] = 1'b0; 
    assign out[9981] = 1'b0; 
    assign out[9982] = 1'b0; 
    assign out[9983] = 1'b0; 
    assign out[9984] = 1'b0; 
    assign out[9985] = 1'b0; 
    assign out[9986] = 1'b0; 
    assign out[9987] = 1'b0; 
    assign out[9988] = 1'b0; 
    assign out[9989] = 1'b0; 
    assign out[9990] = 1'b0; 
    assign out[9991] = 1'b0; 
    assign out[9992] = 1'b0; 
    assign out[9993] = 1'b0; 
    assign out[9994] = 1'b0; 
    assign out[9995] = 1'b0; 
    assign out[9996] = 1'b0; 
    assign out[9997] = 1'b0; 
    assign out[9998] = 1'b0; 
    assign out[9999] = 1'b0; 
    assign out[10000] = 1'b0; 
    assign out[10001] = 1'b0; 
    assign out[10002] = 1'b0; 
    assign out[10003] = 1'b0; 
    assign out[10004] = 1'b0; 
    assign out[10005] = 1'b0; 
    assign out[10006] = 1'b0; 
    assign out[10007] = 1'b0; 
    assign out[10008] = 1'b0; 
    assign out[10009] = 1'b0; 
    assign out[10010] = 1'b0; 
    assign out[10011] = 1'b0; 
    assign out[10012] = 1'b0; 
    assign out[10013] = 1'b0; 
    assign out[10014] = 1'b0; 
    assign out[10015] = 1'b0; 
    assign out[10016] = 1'b0; 
    assign out[10017] = 1'b0; 
    assign out[10018] = 1'b0; 
    assign out[10019] = 1'b0; 
    assign out[10020] = 1'b0; 
    assign out[10021] = 1'b0; 
    assign out[10022] = 1'b0; 
    assign out[10023] = 1'b0; 
    assign out[10024] = 1'b0; 
    assign out[10025] = 1'b0; 
    assign out[10026] = 1'b0; 
    assign out[10027] = 1'b0; 
    assign out[10028] = 1'b0; 
    assign out[10029] = 1'b0; 
    assign out[10030] = 1'b0; 
    assign out[10031] = 1'b0; 
    assign out[10032] = 1'b0; 
    assign out[10033] = 1'b0; 
    assign out[10034] = 1'b0; 
    assign out[10035] = 1'b0; 
    assign out[10036] = 1'b0; 
    assign out[10037] = 1'b0; 
    assign out[10038] = 1'b0; 
    assign out[10039] = 1'b0; 
    assign out[10040] = 1'b0; 
    assign out[10041] = 1'b0; 
    assign out[10042] = 1'b0; 
    assign out[10043] = 1'b0; 
    assign out[10044] = 1'b0; 
    assign out[10045] = 1'b0; 
    assign out[10046] = 1'b0; 
    assign out[10047] = 1'b0; 
    assign out[10048] = 1'b0; 
    assign out[10049] = 1'b0; 
    assign out[10050] = 1'b0; 
    assign out[10051] = 1'b0; 
    assign out[10052] = 1'b0; 
    assign out[10053] = 1'b0; 
    assign out[10054] = 1'b0; 
    assign out[10055] = 1'b0; 
    assign out[10056] = 1'b0; 
    assign out[10057] = 1'b0; 
    assign out[10058] = 1'b0; 
    assign out[10059] = 1'b0; 
    assign out[10060] = 1'b0; 
    assign out[10061] = 1'b0; 
    assign out[10062] = 1'b0; 
    assign out[10063] = 1'b0; 
    assign out[10064] = 1'b0; 
    assign out[10065] = 1'b0; 
    assign out[10066] = 1'b0; 
    assign out[10067] = 1'b0; 
    assign out[10068] = 1'b0; 
    assign out[10069] = 1'b0; 
    assign out[10070] = 1'b0; 
    assign out[10071] = 1'b0; 
    assign out[10072] = 1'b0; 
    assign out[10073] = 1'b0; 
    assign out[10074] = 1'b0; 
    assign out[10075] = 1'b0; 
    assign out[10076] = 1'b0; 
    assign out[10077] = 1'b0; 
    assign out[10078] = 1'b0; 
    assign out[10079] = 1'b0; 
    assign out[10080] = 1'b0; 
    assign out[10081] = 1'b0; 
    assign out[10082] = 1'b0; 
    assign out[10083] = 1'b0; 
    assign out[10084] = 1'b0; 
    assign out[10085] = 1'b0; 
    assign out[10086] = 1'b0; 
    assign out[10087] = 1'b0; 
    assign out[10088] = 1'b0; 
    assign out[10089] = 1'b0; 
    assign out[10090] = 1'b0; 
    assign out[10091] = 1'b0; 
    assign out[10092] = 1'b0; 
    assign out[10093] = 1'b0; 
    assign out[10094] = 1'b0; 
    assign out[10095] = 1'b0; 
    assign out[10096] = 1'b0; 
    assign out[10097] = 1'b0; 
    assign out[10098] = 1'b0; 
    assign out[10099] = 1'b0; 
    assign out[10100] = 1'b0; 
    assign out[10101] = 1'b0; 
    assign out[10102] = 1'b0; 
    assign out[10103] = 1'b0; 
    assign out[10104] = 1'b0; 
    assign out[10105] = 1'b0; 
    assign out[10106] = 1'b0; 
    assign out[10107] = 1'b0; 
    assign out[10108] = 1'b0; 
    assign out[10109] = 1'b0; 
    assign out[10110] = 1'b0; 
    assign out[10111] = 1'b0; 
    assign out[10112] = 1'b0; 
    assign out[10113] = 1'b0; 
    assign out[10114] = 1'b0; 
    assign out[10115] = 1'b0; 
    assign out[10116] = 1'b0; 
    assign out[10117] = 1'b0; 
    assign out[10118] = 1'b0; 
    assign out[10119] = 1'b0; 
    assign out[10120] = 1'b0; 
    assign out[10121] = 1'b0; 
    assign out[10122] = 1'b0; 
    assign out[10123] = 1'b0; 
    assign out[10124] = 1'b0; 
    assign out[10125] = 1'b0; 
    assign out[10126] = 1'b0; 
    assign out[10127] = 1'b0; 
    assign out[10128] = 1'b0; 
    assign out[10129] = 1'b0; 
    assign out[10130] = 1'b0; 
    assign out[10131] = 1'b0; 
    assign out[10132] = 1'b0; 
    assign out[10133] = 1'b0; 
    assign out[10134] = 1'b0; 
    assign out[10135] = 1'b0; 
    assign out[10136] = 1'b0; 
    assign out[10137] = 1'b0; 
    assign out[10138] = 1'b0; 
    assign out[10139] = 1'b0; 
    assign out[10140] = 1'b0; 
    assign out[10141] = 1'b0; 
    assign out[10142] = 1'b0; 
    assign out[10143] = 1'b0; 
    assign out[10144] = 1'b0; 
    assign out[10145] = 1'b0; 
    assign out[10146] = 1'b0; 
    assign out[10147] = 1'b0; 
    assign out[10148] = 1'b0; 
    assign out[10149] = 1'b0; 
    assign out[10150] = 1'b0; 
    assign out[10151] = 1'b0; 
    assign out[10152] = 1'b0; 
    assign out[10153] = 1'b0; 
    assign out[10154] = 1'b0; 
    assign out[10155] = 1'b0; 
    assign out[10156] = 1'b0; 
    assign out[10157] = 1'b0; 
    assign out[10158] = 1'b0; 
    assign out[10159] = 1'b0; 
    assign out[10160] = 1'b0; 
    assign out[10161] = 1'b0; 
    assign out[10162] = 1'b0; 
    assign out[10163] = 1'b0; 
    assign out[10164] = 1'b0; 
    assign out[10165] = 1'b0; 
    assign out[10166] = 1'b0; 
    assign out[10167] = 1'b0; 
    assign out[10168] = 1'b0; 
    assign out[10169] = 1'b0; 
    assign out[10170] = 1'b0; 
    assign out[10171] = 1'b0; 
    assign out[10172] = 1'b0; 
    assign out[10173] = 1'b0; 
    assign out[10174] = 1'b0; 
    assign out[10175] = 1'b0; 
    assign out[10176] = 1'b0; 
    assign out[10177] = 1'b0; 
    assign out[10178] = 1'b0; 
    assign out[10179] = 1'b0; 
    assign out[10180] = 1'b0; 
    assign out[10181] = 1'b0; 
    assign out[10182] = 1'b0; 
    assign out[10183] = 1'b0; 
    assign out[10184] = 1'b0; 
    assign out[10185] = 1'b0; 
    assign out[10186] = 1'b0; 
    assign out[10187] = 1'b0; 
    assign out[10188] = 1'b0; 
    assign out[10189] = 1'b0; 
    assign out[10190] = 1'b0; 
    assign out[10191] = 1'b0; 
    assign out[10192] = 1'b0; 
    assign out[10193] = 1'b0; 
    assign out[10194] = 1'b0; 
    assign out[10195] = 1'b0; 
    assign out[10196] = 1'b0; 
    assign out[10197] = 1'b0; 
    assign out[10198] = 1'b0; 
    assign out[10199] = 1'b0; 
    assign out[10200] = 1'b0; 
    assign out[10201] = 1'b0; 
    assign out[10202] = 1'b0; 
    assign out[10203] = 1'b0; 
    assign out[10204] = 1'b0; 
    assign out[10205] = 1'b0; 
    assign out[10206] = 1'b0; 
    assign out[10207] = 1'b0; 
    assign out[10208] = 1'b0; 
    assign out[10209] = 1'b0; 
    assign out[10210] = 1'b0; 
    assign out[10211] = 1'b0; 
    assign out[10212] = 1'b0; 
    assign out[10213] = 1'b0; 
    assign out[10214] = 1'b0; 
    assign out[10215] = 1'b0; 
    assign out[10216] = 1'b0; 
    assign out[10217] = 1'b0; 
    assign out[10218] = 1'b0; 
    assign out[10219] = 1'b0; 
    assign out[10220] = 1'b0; 
    assign out[10221] = 1'b0; 
    assign out[10222] = 1'b0; 
    assign out[10223] = 1'b0; 
    assign out[10224] = 1'b0; 
    assign out[10225] = 1'b0; 
    assign out[10226] = 1'b0; 
    assign out[10227] = 1'b0; 
    assign out[10228] = 1'b0; 
    assign out[10229] = 1'b0; 
    assign out[10230] = 1'b0; 
    assign out[10231] = 1'b0; 
    assign out[10232] = 1'b0; 
    assign out[10233] = 1'b0; 
    assign out[10234] = 1'b0; 
    assign out[10235] = 1'b0; 
    assign out[10236] = 1'b0; 
    assign out[10237] = 1'b0; 
    assign out[10238] = 1'b0; 
    assign out[10239] = 1'b0; 
    assign out[10240] = 1'b0; 
    assign out[10241] = 1'b0; 
    assign out[10242] = 1'b0; 
    assign out[10243] = 1'b0; 
    assign out[10244] = 1'b0; 
    assign out[10245] = 1'b0; 
    assign out[10246] = 1'b0; 
    assign out[10247] = 1'b0; 
    assign out[10248] = 1'b0; 
    assign out[10249] = 1'b0; 
    assign out[10250] = 1'b0; 
    assign out[10251] = 1'b0; 
    assign out[10252] = 1'b0; 
    assign out[10253] = 1'b0; 
    assign out[10254] = 1'b0; 
    assign out[10255] = 1'b0; 
    assign out[10256] = 1'b0; 
    assign out[10257] = 1'b0; 
    assign out[10258] = 1'b0; 
    assign out[10259] = 1'b0; 
    assign out[10260] = 1'b0; 
    assign out[10261] = 1'b0; 
    assign out[10262] = 1'b0; 
    assign out[10263] = 1'b0; 
    assign out[10264] = 1'b0; 
    assign out[10265] = 1'b0; 
    assign out[10266] = 1'b0; 
    assign out[10267] = 1'b0; 
    assign out[10268] = 1'b0; 
    assign out[10269] = 1'b0; 
    assign out[10270] = 1'b0; 
    assign out[10271] = 1'b0; 
    assign out[10272] = 1'b0; 
    assign out[10273] = 1'b0; 
    assign out[10274] = 1'b0; 
    assign out[10275] = 1'b0; 
    assign out[10276] = 1'b0; 
    assign out[10277] = 1'b0; 
    assign out[10278] = 1'b0; 
    assign out[10279] = 1'b0; 
    assign out[10280] = 1'b0; 
    assign out[10281] = 1'b0; 
    assign out[10282] = 1'b0; 
    assign out[10283] = 1'b0; 
    assign out[10284] = 1'b0; 
    assign out[10285] = 1'b0; 
    assign out[10286] = 1'b0; 
    assign out[10287] = 1'b0; 
    assign out[10288] = 1'b0; 
    assign out[10289] = 1'b0; 
    assign out[10290] = 1'b0; 
    assign out[10291] = 1'b0; 
    assign out[10292] = 1'b0; 
    assign out[10293] = 1'b0; 
    assign out[10294] = 1'b0; 
    assign out[10295] = 1'b0; 
    assign out[10296] = 1'b0; 
    assign out[10297] = 1'b0; 
    assign out[10298] = 1'b0; 
    assign out[10299] = 1'b0; 
    assign out[10300] = 1'b0; 
    assign out[10301] = 1'b0; 
    assign out[10302] = 1'b0; 
    assign out[10303] = 1'b0; 
    assign out[10304] = 1'b0; 
    assign out[10305] = 1'b0; 
    assign out[10306] = 1'b0; 
    assign out[10307] = 1'b0; 
    assign out[10308] = 1'b0; 
    assign out[10309] = 1'b0; 
    assign out[10310] = 1'b0; 
    assign out[10311] = 1'b0; 
    assign out[10312] = 1'b0; 
    assign out[10313] = 1'b0; 
    assign out[10314] = 1'b0; 
    assign out[10315] = 1'b0; 
    assign out[10316] = 1'b0; 
    assign out[10317] = 1'b0; 
    assign out[10318] = 1'b0; 
    assign out[10319] = 1'b0; 
    assign out[10320] = 1'b0; 
    assign out[10321] = 1'b0; 
    assign out[10322] = 1'b0; 
    assign out[10323] = 1'b0; 
    assign out[10324] = 1'b0; 
    assign out[10325] = 1'b0; 
    assign out[10326] = 1'b0; 
    assign out[10327] = 1'b0; 
    assign out[10328] = 1'b0; 
    assign out[10329] = 1'b0; 
    assign out[10330] = 1'b0; 
    assign out[10331] = 1'b0; 
    assign out[10332] = 1'b0; 
    assign out[10333] = 1'b0; 
    assign out[10334] = 1'b0; 
    assign out[10335] = 1'b0; 
    assign out[10336] = 1'b0; 
    assign out[10337] = 1'b0; 
    assign out[10338] = 1'b0; 
    assign out[10339] = 1'b0; 
    assign out[10340] = 1'b0; 
    assign out[10341] = 1'b0; 
    assign out[10342] = 1'b0; 
    assign out[10343] = 1'b0; 
    assign out[10344] = 1'b0; 
    assign out[10345] = 1'b0; 
    assign out[10346] = 1'b0; 
    assign out[10347] = 1'b0; 
    assign out[10348] = 1'b0; 
    assign out[10349] = 1'b0; 
    assign out[10350] = 1'b0; 
    assign out[10351] = 1'b0; 
    assign out[10352] = 1'b0; 
    assign out[10353] = 1'b0; 
    assign out[10354] = 1'b0; 
    assign out[10355] = 1'b0; 
    assign out[10356] = 1'b0; 
    assign out[10357] = 1'b0; 
    assign out[10358] = 1'b0; 
    assign out[10359] = 1'b0; 
    assign out[10360] = 1'b0; 
    assign out[10361] = 1'b0; 
    assign out[10362] = 1'b0; 
    assign out[10363] = 1'b0; 
    assign out[10364] = 1'b0; 
    assign out[10365] = 1'b0; 
    assign out[10366] = 1'b0; 
    assign out[10367] = 1'b0; 
    assign out[10368] = 1'b0; 
    assign out[10369] = 1'b0; 
    assign out[10370] = 1'b0; 
    assign out[10371] = 1'b0; 
    assign out[10372] = 1'b0; 
    assign out[10373] = 1'b0; 
    assign out[10374] = 1'b0; 
    assign out[10375] = 1'b0; 
    assign out[10376] = 1'b0; 
    assign out[10377] = 1'b0; 
    assign out[10378] = 1'b0; 
    assign out[10379] = 1'b0; 
    assign out[10380] = 1'b0; 
    assign out[10381] = 1'b0; 
    assign out[10382] = 1'b0; 
    assign out[10383] = 1'b0; 
    assign out[10384] = 1'b0; 
    assign out[10385] = 1'b0; 
    assign out[10386] = 1'b0; 
    assign out[10387] = 1'b0; 
    assign out[10388] = 1'b0; 
    assign out[10389] = 1'b0; 
    assign out[10390] = 1'b0; 
    assign out[10391] = 1'b0; 
    assign out[10392] = 1'b0; 
    assign out[10393] = 1'b0; 
    assign out[10394] = 1'b0; 
    assign out[10395] = 1'b0; 
    assign out[10396] = 1'b0; 
    assign out[10397] = 1'b0; 
    assign out[10398] = 1'b0; 
    assign out[10399] = 1'b0; 
    assign out[10400] = 1'b0; 
    assign out[10401] = 1'b0; 
    assign out[10402] = 1'b0; 
    assign out[10403] = 1'b0; 
    assign out[10404] = 1'b0; 
    assign out[10405] = 1'b0; 
    assign out[10406] = 1'b0; 
    assign out[10407] = 1'b0; 
    assign out[10408] = 1'b0; 
    assign out[10409] = 1'b0; 
    assign out[10410] = 1'b0; 
    assign out[10411] = 1'b0; 
    assign out[10412] = 1'b0; 
    assign out[10413] = 1'b0; 
    assign out[10414] = 1'b0; 
    assign out[10415] = 1'b0; 
    assign out[10416] = 1'b0; 
    assign out[10417] = 1'b0; 
    assign out[10418] = 1'b0; 
    assign out[10419] = 1'b0; 
    assign out[10420] = 1'b0; 
    assign out[10421] = 1'b0; 
    assign out[10422] = 1'b0; 
    assign out[10423] = 1'b0; 
    assign out[10424] = 1'b0; 
    assign out[10425] = 1'b0; 
    assign out[10426] = 1'b0; 
    assign out[10427] = 1'b0; 
    assign out[10428] = 1'b0; 
    assign out[10429] = 1'b0; 
    assign out[10430] = 1'b0; 
    assign out[10431] = 1'b0; 
    assign out[10432] = 1'b0; 
    assign out[10433] = 1'b0; 
    assign out[10434] = 1'b0; 
    assign out[10435] = 1'b0; 
    assign out[10436] = 1'b0; 
    assign out[10437] = 1'b0; 
    assign out[10438] = 1'b0; 
    assign out[10439] = 1'b0; 
    assign out[10440] = 1'b0; 
    assign out[10441] = 1'b0; 
    assign out[10442] = 1'b0; 
    assign out[10443] = 1'b0; 
    assign out[10444] = 1'b0; 
    assign out[10445] = 1'b0; 
    assign out[10446] = 1'b0; 
    assign out[10447] = 1'b0; 
    assign out[10448] = 1'b0; 
    assign out[10449] = 1'b0; 
    assign out[10450] = 1'b0; 
    assign out[10451] = 1'b0; 
    assign out[10452] = 1'b0; 
    assign out[10453] = 1'b0; 
    assign out[10454] = 1'b0; 
    assign out[10455] = 1'b0; 
    assign out[10456] = 1'b0; 
    assign out[10457] = 1'b0; 
    assign out[10458] = 1'b0; 
    assign out[10459] = 1'b0; 
    assign out[10460] = 1'b0; 
    assign out[10461] = 1'b0; 
    assign out[10462] = 1'b0; 
    assign out[10463] = 1'b0; 
    assign out[10464] = 1'b0; 
    assign out[10465] = 1'b0; 
    assign out[10466] = 1'b0; 
    assign out[10467] = 1'b0; 
    assign out[10468] = 1'b0; 
    assign out[10469] = 1'b0; 
    assign out[10470] = 1'b0; 
    assign out[10471] = 1'b0; 
    assign out[10472] = 1'b0; 
    assign out[10473] = 1'b0; 
    assign out[10474] = 1'b0; 
    assign out[10475] = 1'b0; 
    assign out[10476] = 1'b0; 
    assign out[10477] = 1'b0; 
    assign out[10478] = 1'b0; 
    assign out[10479] = 1'b0; 
    assign out[10480] = 1'b0; 
    assign out[10481] = 1'b0; 
    assign out[10482] = 1'b0; 
    assign out[10483] = 1'b0; 
    assign out[10484] = 1'b0; 
    assign out[10485] = 1'b0; 
    assign out[10486] = 1'b0; 
    assign out[10487] = 1'b0; 
    assign out[10488] = 1'b0; 
    assign out[10489] = 1'b0; 
    assign out[10490] = 1'b0; 
    assign out[10491] = 1'b0; 
    assign out[10492] = 1'b0; 
    assign out[10493] = 1'b0; 
    assign out[10494] = 1'b0; 
    assign out[10495] = 1'b0; 
    assign out[10496] = 1'b0; 
    assign out[10497] = 1'b0; 
    assign out[10498] = 1'b0; 
    assign out[10499] = 1'b0; 
    assign out[10500] = 1'b0; 
    assign out[10501] = 1'b0; 
    assign out[10502] = 1'b0; 
    assign out[10503] = 1'b0; 
    assign out[10504] = 1'b0; 
    assign out[10505] = 1'b0; 
    assign out[10506] = 1'b0; 
    assign out[10507] = 1'b0; 
    assign out[10508] = 1'b0; 
    assign out[10509] = 1'b0; 
    assign out[10510] = 1'b0; 
    assign out[10511] = 1'b0; 
    assign out[10512] = 1'b0; 
    assign out[10513] = 1'b0; 
    assign out[10514] = 1'b0; 
    assign out[10515] = 1'b0; 
    assign out[10516] = 1'b0; 
    assign out[10517] = 1'b0; 
    assign out[10518] = 1'b0; 
    assign out[10519] = 1'b0; 
    assign out[10520] = 1'b0; 
    assign out[10521] = 1'b0; 
    assign out[10522] = 1'b0; 
    assign out[10523] = 1'b0; 
    assign out[10524] = 1'b0; 
    assign out[10525] = 1'b0; 
    assign out[10526] = 1'b0; 
    assign out[10527] = 1'b0; 
    assign out[10528] = 1'b0; 
    assign out[10529] = 1'b0; 
    assign out[10530] = 1'b0; 
    assign out[10531] = 1'b0; 
    assign out[10532] = 1'b0; 
    assign out[10533] = 1'b0; 
    assign out[10534] = 1'b0; 
    assign out[10535] = 1'b0; 
    assign out[10536] = 1'b0; 
    assign out[10537] = 1'b0; 
    assign out[10538] = 1'b0; 
    assign out[10539] = 1'b0; 
    assign out[10540] = 1'b0; 
    assign out[10541] = 1'b0; 
    assign out[10542] = 1'b0; 
    assign out[10543] = 1'b0; 
    assign out[10544] = 1'b0; 
    assign out[10545] = 1'b0; 
    assign out[10546] = 1'b0; 
    assign out[10547] = 1'b0; 
    assign out[10548] = 1'b0; 
    assign out[10549] = 1'b0; 
    assign out[10550] = 1'b0; 
    assign out[10551] = 1'b0; 
    assign out[10552] = 1'b0; 
    assign out[10553] = 1'b0; 
    assign out[10554] = 1'b0; 
    assign out[10555] = 1'b0; 
    assign out[10556] = 1'b0; 
    assign out[10557] = 1'b0; 
    assign out[10558] = 1'b0; 
    assign out[10559] = 1'b0; 
    assign out[10560] = 1'b0; 
    assign out[10561] = 1'b0; 
    assign out[10562] = 1'b0; 
    assign out[10563] = 1'b0; 
    assign out[10564] = 1'b0; 
    assign out[10565] = 1'b0; 
    assign out[10566] = 1'b0; 
    assign out[10567] = 1'b0; 
    assign out[10568] = 1'b0; 
    assign out[10569] = 1'b0; 
    assign out[10570] = 1'b0; 
    assign out[10571] = 1'b0; 
    assign out[10572] = 1'b0; 
    assign out[10573] = 1'b0; 
    assign out[10574] = 1'b0; 
    assign out[10575] = 1'b0; 
    assign out[10576] = 1'b0; 
    assign out[10577] = 1'b0; 
    assign out[10578] = 1'b0; 
    assign out[10579] = 1'b0; 
    assign out[10580] = 1'b0; 
    assign out[10581] = 1'b0; 
    assign out[10582] = 1'b0; 
    assign out[10583] = 1'b0; 
    assign out[10584] = 1'b0; 
    assign out[10585] = 1'b0; 
    assign out[10586] = 1'b0; 
    assign out[10587] = 1'b0; 
    assign out[10588] = 1'b0; 
    assign out[10589] = 1'b0; 
    assign out[10590] = 1'b0; 
    assign out[10591] = 1'b0; 
    assign out[10592] = 1'b0; 
    assign out[10593] = 1'b0; 
    assign out[10594] = 1'b0; 
    assign out[10595] = 1'b0; 
    assign out[10596] = 1'b0; 
    assign out[10597] = 1'b0; 
    assign out[10598] = 1'b0; 
    assign out[10599] = 1'b0; 
    assign out[10600] = 1'b0; 
    assign out[10601] = 1'b0; 
    assign out[10602] = 1'b0; 
    assign out[10603] = 1'b0; 
    assign out[10604] = 1'b0; 
    assign out[10605] = 1'b0; 
    assign out[10606] = 1'b0; 
    assign out[10607] = 1'b0; 
    assign out[10608] = 1'b0; 
    assign out[10609] = 1'b0; 
    assign out[10610] = 1'b0; 
    assign out[10611] = 1'b0; 
    assign out[10612] = 1'b0; 
    assign out[10613] = 1'b0; 
    assign out[10614] = 1'b0; 
    assign out[10615] = 1'b0; 
    assign out[10616] = 1'b0; 
    assign out[10617] = 1'b0; 
    assign out[10618] = 1'b0; 
    assign out[10619] = 1'b0; 
    assign out[10620] = 1'b0; 
    assign out[10621] = 1'b0; 
    assign out[10622] = 1'b0; 
    assign out[10623] = 1'b0; 
    assign out[10624] = 1'b0; 
    assign out[10625] = 1'b0; 
    assign out[10626] = 1'b0; 
    assign out[10627] = 1'b0; 
    assign out[10628] = 1'b0; 
    assign out[10629] = 1'b0; 
    assign out[10630] = 1'b0; 
    assign out[10631] = 1'b0; 
    assign out[10632] = 1'b0; 
    assign out[10633] = 1'b0; 
    assign out[10634] = 1'b0; 
    assign out[10635] = 1'b0; 
    assign out[10636] = 1'b0; 
    assign out[10637] = 1'b0; 
    assign out[10638] = 1'b0; 
    assign out[10639] = 1'b0; 
    assign out[10640] = 1'b0; 
    assign out[10641] = 1'b0; 
    assign out[10642] = 1'b0; 
    assign out[10643] = 1'b0; 
    assign out[10644] = 1'b0; 
    assign out[10645] = 1'b0; 
    assign out[10646] = 1'b0; 
    assign out[10647] = 1'b0; 
    assign out[10648] = 1'b0; 
    assign out[10649] = 1'b0; 
    assign out[10650] = 1'b0; 
    assign out[10651] = 1'b0; 
    assign out[10652] = 1'b0; 
    assign out[10653] = 1'b0; 
    assign out[10654] = 1'b0; 
    assign out[10655] = 1'b0; 
    assign out[10656] = 1'b0; 
    assign out[10657] = 1'b0; 
    assign out[10658] = 1'b0; 
    assign out[10659] = 1'b0; 
    assign out[10660] = 1'b0; 
    assign out[10661] = 1'b0; 
    assign out[10662] = 1'b0; 
    assign out[10663] = 1'b0; 
    assign out[10664] = 1'b0; 
    assign out[10665] = 1'b0; 
    assign out[10666] = 1'b0; 
    assign out[10667] = 1'b0; 
    assign out[10668] = 1'b0; 
    assign out[10669] = 1'b0; 
    assign out[10670] = 1'b0; 
    assign out[10671] = 1'b0; 
    assign out[10672] = 1'b0; 
    assign out[10673] = 1'b0; 
    assign out[10674] = 1'b0; 
    assign out[10675] = 1'b0; 
    assign out[10676] = 1'b0; 
    assign out[10677] = 1'b0; 
    assign out[10678] = 1'b0; 
    assign out[10679] = 1'b0; 
    assign out[10680] = 1'b0; 
    assign out[10681] = 1'b0; 
    assign out[10682] = 1'b0; 
    assign out[10683] = 1'b0; 
    assign out[10684] = 1'b0; 
    assign out[10685] = 1'b0; 
    assign out[10686] = 1'b0; 
    assign out[10687] = 1'b0; 
    assign out[10688] = 1'b0; 
    assign out[10689] = 1'b0; 
    assign out[10690] = 1'b0; 
    assign out[10691] = 1'b0; 
    assign out[10692] = 1'b0; 
    assign out[10693] = 1'b0; 
    assign out[10694] = 1'b0; 
    assign out[10695] = 1'b0; 
    assign out[10696] = 1'b0; 
    assign out[10697] = 1'b0; 
    assign out[10698] = 1'b0; 
    assign out[10699] = 1'b0; 
    assign out[10700] = 1'b0; 
    assign out[10701] = 1'b0; 
    assign out[10702] = 1'b0; 
    assign out[10703] = 1'b0; 
    assign out[10704] = 1'b0; 
    assign out[10705] = 1'b0; 
    assign out[10706] = 1'b0; 
    assign out[10707] = 1'b0; 
    assign out[10708] = 1'b0; 
    assign out[10709] = 1'b0; 
    assign out[10710] = 1'b0; 
    assign out[10711] = 1'b0; 
    assign out[10712] = 1'b0; 
    assign out[10713] = 1'b0; 
    assign out[10714] = 1'b0; 
    assign out[10715] = 1'b0; 
    assign out[10716] = 1'b0; 
    assign out[10717] = 1'b0; 
    assign out[10718] = 1'b0; 
    assign out[10719] = 1'b0; 
    assign out[10720] = 1'b0; 
    assign out[10721] = 1'b0; 
    assign out[10722] = 1'b0; 
    assign out[10723] = 1'b0; 
    assign out[10724] = 1'b0; 
    assign out[10725] = 1'b0; 
    assign out[10726] = 1'b0; 
    assign out[10727] = 1'b0; 
    assign out[10728] = 1'b0; 
    assign out[10729] = 1'b0; 
    assign out[10730] = 1'b0; 
    assign out[10731] = 1'b0; 
    assign out[10732] = 1'b0; 
    assign out[10733] = 1'b0; 
    assign out[10734] = 1'b0; 
    assign out[10735] = 1'b0; 
    assign out[10736] = 1'b0; 
    assign out[10737] = 1'b0; 
    assign out[10738] = 1'b0; 
    assign out[10739] = 1'b0; 
    assign out[10740] = 1'b0; 
    assign out[10741] = 1'b0; 
    assign out[10742] = 1'b0; 
    assign out[10743] = 1'b0; 
    assign out[10744] = 1'b0; 
    assign out[10745] = 1'b0; 
    assign out[10746] = 1'b0; 
    assign out[10747] = 1'b0; 
    assign out[10748] = 1'b0; 
    assign out[10749] = 1'b0; 
    assign out[10750] = 1'b0; 
    assign out[10751] = 1'b0; 
    assign out[10752] = 1'b0; 
    assign out[10753] = 1'b0; 
    assign out[10754] = 1'b0; 
    assign out[10755] = 1'b0; 
    assign out[10756] = 1'b0; 
    assign out[10757] = 1'b0; 
    assign out[10758] = 1'b0; 
    assign out[10759] = 1'b0; 
    assign out[10760] = 1'b0; 
    assign out[10761] = 1'b0; 
    assign out[10762] = 1'b0; 
    assign out[10763] = 1'b0; 
    assign out[10764] = 1'b0; 
    assign out[10765] = 1'b0; 
    assign out[10766] = 1'b0; 
    assign out[10767] = 1'b0; 
    assign out[10768] = 1'b0; 
    assign out[10769] = 1'b0; 
    assign out[10770] = 1'b0; 
    assign out[10771] = 1'b0; 
    assign out[10772] = 1'b0; 
    assign out[10773] = 1'b0; 
    assign out[10774] = 1'b0; 
    assign out[10775] = 1'b0; 
    assign out[10776] = 1'b0; 
    assign out[10777] = 1'b0; 
    assign out[10778] = 1'b0; 
    assign out[10779] = 1'b0; 
    assign out[10780] = 1'b0; 
    assign out[10781] = 1'b0; 
    assign out[10782] = 1'b0; 
    assign out[10783] = 1'b0; 
    assign out[10784] = 1'b0; 
    assign out[10785] = 1'b0; 
    assign out[10786] = 1'b0; 
    assign out[10787] = 1'b0; 
    assign out[10788] = 1'b0; 
    assign out[10789] = 1'b0; 
    assign out[10790] = 1'b0; 
    assign out[10791] = 1'b0; 
    assign out[10792] = 1'b0; 
    assign out[10793] = 1'b0; 
    assign out[10794] = 1'b0; 
    assign out[10795] = 1'b0; 
    assign out[10796] = 1'b0; 
    assign out[10797] = 1'b0; 
    assign out[10798] = 1'b0; 
    assign out[10799] = 1'b0; 
    assign out[10800] = 1'b0; 
    assign out[10801] = 1'b0; 
    assign out[10802] = 1'b0; 
    assign out[10803] = 1'b0; 
    assign out[10804] = 1'b0; 
    assign out[10805] = 1'b0; 
    assign out[10806] = 1'b0; 
    assign out[10807] = 1'b0; 
    assign out[10808] = 1'b0; 
    assign out[10809] = 1'b0; 
    assign out[10810] = 1'b0; 
    assign out[10811] = 1'b0; 
    assign out[10812] = 1'b0; 
    assign out[10813] = 1'b0; 
    assign out[10814] = 1'b0; 
    assign out[10815] = 1'b0; 
    assign out[10816] = 1'b0; 
    assign out[10817] = 1'b0; 
    assign out[10818] = 1'b0; 
    assign out[10819] = 1'b0; 
    assign out[10820] = 1'b0; 
    assign out[10821] = 1'b0; 
    assign out[10822] = 1'b0; 
    assign out[10823] = 1'b0; 
    assign out[10824] = 1'b0; 
    assign out[10825] = 1'b0; 
    assign out[10826] = 1'b0; 
    assign out[10827] = 1'b0; 
    assign out[10828] = 1'b0; 
    assign out[10829] = 1'b0; 
    assign out[10830] = 1'b0; 
    assign out[10831] = 1'b0; 
    assign out[10832] = 1'b0; 
    assign out[10833] = 1'b0; 
    assign out[10834] = 1'b0; 
    assign out[10835] = 1'b0; 
    assign out[10836] = 1'b0; 
    assign out[10837] = 1'b0; 
    assign out[10838] = 1'b0; 
    assign out[10839] = 1'b0; 
    assign out[10840] = 1'b0; 
    assign out[10841] = 1'b0; 
    assign out[10842] = 1'b0; 
    assign out[10843] = 1'b0; 
    assign out[10844] = 1'b0; 
    assign out[10845] = 1'b0; 
    assign out[10846] = 1'b0; 
    assign out[10847] = 1'b0; 
    assign out[10848] = 1'b0; 
    assign out[10849] = 1'b0; 
    assign out[10850] = 1'b0; 
    assign out[10851] = 1'b0; 
    assign out[10852] = 1'b0; 
    assign out[10853] = 1'b0; 
    assign out[10854] = 1'b0; 
    assign out[10855] = 1'b0; 
    assign out[10856] = 1'b0; 
    assign out[10857] = 1'b0; 
    assign out[10858] = 1'b0; 
    assign out[10859] = 1'b0; 
    assign out[10860] = 1'b0; 
    assign out[10861] = 1'b0; 
    assign out[10862] = 1'b0; 
    assign out[10863] = 1'b0; 
    assign out[10864] = 1'b0; 
    assign out[10865] = 1'b0; 
    assign out[10866] = 1'b0; 
    assign out[10867] = 1'b0; 
    assign out[10868] = 1'b0; 
    assign out[10869] = 1'b0; 
    assign out[10870] = 1'b0; 
    assign out[10871] = 1'b0; 
    assign out[10872] = 1'b0; 
    assign out[10873] = 1'b0; 
    assign out[10874] = 1'b0; 
    assign out[10875] = 1'b0; 
    assign out[10876] = 1'b0; 
    assign out[10877] = 1'b0; 
    assign out[10878] = 1'b0; 
    assign out[10879] = 1'b0; 
    assign out[10880] = 1'b0; 
    assign out[10881] = 1'b0; 
    assign out[10882] = 1'b0; 
    assign out[10883] = 1'b0; 
    assign out[10884] = 1'b0; 
    assign out[10885] = 1'b0; 
    assign out[10886] = 1'b0; 
    assign out[10887] = 1'b0; 
    assign out[10888] = 1'b0; 
    assign out[10889] = 1'b0; 
    assign out[10890] = 1'b0; 
    assign out[10891] = 1'b0; 
    assign out[10892] = 1'b0; 
    assign out[10893] = 1'b0; 
    assign out[10894] = 1'b0; 
    assign out[10895] = 1'b0; 
    assign out[10896] = 1'b0; 
    assign out[10897] = 1'b0; 
    assign out[10898] = 1'b0; 
    assign out[10899] = 1'b0; 
    assign out[10900] = 1'b0; 
    assign out[10901] = 1'b0; 
    assign out[10902] = 1'b0; 
    assign out[10903] = 1'b0; 
    assign out[10904] = 1'b0; 
    assign out[10905] = 1'b0; 
    assign out[10906] = 1'b0; 
    assign out[10907] = 1'b0; 
    assign out[10908] = 1'b0; 
    assign out[10909] = 1'b0; 
    assign out[10910] = 1'b0; 
    assign out[10911] = 1'b0; 
    assign out[10912] = 1'b0; 
    assign out[10913] = 1'b0; 
    assign out[10914] = 1'b0; 
    assign out[10915] = 1'b0; 
    assign out[10916] = 1'b0; 
    assign out[10917] = 1'b0; 
    assign out[10918] = 1'b0; 
    assign out[10919] = 1'b0; 
    assign out[10920] = 1'b0; 
    assign out[10921] = 1'b0; 
    assign out[10922] = 1'b0; 
    assign out[10923] = 1'b0; 
    assign out[10924] = 1'b0; 
    assign out[10925] = 1'b0; 
    assign out[10926] = 1'b0; 
    assign out[10927] = 1'b0; 
    assign out[10928] = 1'b0; 
    assign out[10929] = 1'b0; 
    assign out[10930] = 1'b0; 
    assign out[10931] = 1'b0; 
    assign out[10932] = 1'b0; 
    assign out[10933] = 1'b0; 
    assign out[10934] = 1'b0; 
    assign out[10935] = 1'b0; 
    assign out[10936] = 1'b0; 
    assign out[10937] = 1'b0; 
    assign out[10938] = 1'b0; 
    assign out[10939] = 1'b0; 
    assign out[10940] = 1'b0; 
    assign out[10941] = 1'b0; 
    assign out[10942] = 1'b0; 
    assign out[10943] = 1'b0; 
    assign out[10944] = 1'b0; 
    assign out[10945] = 1'b0; 
    assign out[10946] = 1'b0; 
    assign out[10947] = 1'b0; 
    assign out[10948] = 1'b0; 
    assign out[10949] = 1'b0; 
    assign out[10950] = 1'b0; 
    assign out[10951] = 1'b0; 
    assign out[10952] = 1'b0; 
    assign out[10953] = 1'b0; 
    assign out[10954] = 1'b0; 
    assign out[10955] = 1'b0; 
    assign out[10956] = 1'b0; 
    assign out[10957] = 1'b0; 
    assign out[10958] = 1'b0; 
    assign out[10959] = 1'b0; 
    assign out[10960] = 1'b0; 
    assign out[10961] = 1'b0; 
    assign out[10962] = 1'b0; 
    assign out[10963] = 1'b0; 
    assign out[10964] = 1'b0; 
    assign out[10965] = 1'b0; 
    assign out[10966] = 1'b0; 
    assign out[10967] = 1'b0; 
    assign out[10968] = 1'b0; 
    assign out[10969] = 1'b0; 
    assign out[10970] = 1'b0; 
    assign out[10971] = 1'b0; 
    assign out[10972] = 1'b0; 
    assign out[10973] = 1'b0; 
    assign out[10974] = 1'b0; 
    assign out[10975] = 1'b0; 
    assign out[10976] = 1'b0; 
    assign out[10977] = 1'b0; 
    assign out[10978] = 1'b0; 
    assign out[10979] = 1'b0; 
    assign out[10980] = 1'b0; 
    assign out[10981] = 1'b0; 
    assign out[10982] = 1'b0; 
    assign out[10983] = 1'b0; 
    assign out[10984] = 1'b0; 
    assign out[10985] = 1'b0; 
    assign out[10986] = 1'b0; 
    assign out[10987] = 1'b0; 
    assign out[10988] = 1'b0; 
    assign out[10989] = 1'b0; 
    assign out[10990] = 1'b0; 
    assign out[10991] = 1'b0; 
    assign out[10992] = 1'b0; 
    assign out[10993] = 1'b0; 
    assign out[10994] = 1'b0; 
    assign out[10995] = 1'b0; 
    assign out[10996] = 1'b0; 
    assign out[10997] = 1'b0; 
    assign out[10998] = 1'b0; 
    assign out[10999] = 1'b0; 
    assign out[11000] = 1'b0; 
    assign out[11001] = 1'b0; 
    assign out[11002] = 1'b0; 
    assign out[11003] = 1'b0; 
    assign out[11004] = 1'b0; 
    assign out[11005] = 1'b0; 
    assign out[11006] = 1'b0; 
    assign out[11007] = 1'b0; 
    assign out[11008] = 1'b0; 
    assign out[11009] = 1'b0; 
    assign out[11010] = 1'b0; 
    assign out[11011] = 1'b0; 
    assign out[11012] = 1'b0; 
    assign out[11013] = 1'b0; 
    assign out[11014] = 1'b0; 
    assign out[11015] = 1'b0; 
    assign out[11016] = 1'b0; 
    assign out[11017] = 1'b0; 
    assign out[11018] = 1'b0; 
    assign out[11019] = 1'b0; 
    assign out[11020] = 1'b0; 
    assign out[11021] = 1'b0; 
    assign out[11022] = 1'b0; 
    assign out[11023] = 1'b0; 
    assign out[11024] = 1'b0; 
    assign out[11025] = 1'b0; 
    assign out[11026] = 1'b0; 
    assign out[11027] = 1'b0; 
    assign out[11028] = 1'b0; 
    assign out[11029] = 1'b0; 
    assign out[11030] = 1'b0; 
    assign out[11031] = 1'b0; 
    assign out[11032] = 1'b0; 
    assign out[11033] = 1'b0; 
    assign out[11034] = 1'b0; 
    assign out[11035] = 1'b0; 
    assign out[11036] = 1'b0; 
    assign out[11037] = 1'b0; 
    assign out[11038] = 1'b0; 
    assign out[11039] = 1'b0; 
    assign out[11040] = 1'b0; 
    assign out[11041] = 1'b0; 
    assign out[11042] = 1'b0; 
    assign out[11043] = 1'b0; 
    assign out[11044] = 1'b0; 
    assign out[11045] = 1'b0; 
    assign out[11046] = 1'b0; 
    assign out[11047] = 1'b0; 
    assign out[11048] = 1'b0; 
    assign out[11049] = 1'b0; 
    assign out[11050] = 1'b0; 
    assign out[11051] = 1'b0; 
    assign out[11052] = 1'b0; 
    assign out[11053] = 1'b0; 
    assign out[11054] = 1'b0; 
    assign out[11055] = 1'b0; 
    assign out[11056] = 1'b0; 
    assign out[11057] = 1'b0; 
    assign out[11058] = 1'b0; 
    assign out[11059] = 1'b0; 
    assign out[11060] = 1'b0; 
    assign out[11061] = 1'b0; 
    assign out[11062] = 1'b0; 
    assign out[11063] = 1'b0; 
    assign out[11064] = 1'b0; 
    assign out[11065] = 1'b0; 
    assign out[11066] = 1'b0; 
    assign out[11067] = 1'b0; 
    assign out[11068] = 1'b0; 
    assign out[11069] = 1'b0; 
    assign out[11070] = 1'b0; 
    assign out[11071] = 1'b0; 
    assign out[11072] = 1'b0; 
    assign out[11073] = 1'b0; 
    assign out[11074] = 1'b0; 
    assign out[11075] = 1'b0; 
    assign out[11076] = 1'b0; 
    assign out[11077] = 1'b0; 
    assign out[11078] = 1'b0; 
    assign out[11079] = 1'b0; 
    assign out[11080] = 1'b0; 
    assign out[11081] = 1'b0; 
    assign out[11082] = 1'b0; 
    assign out[11083] = 1'b0; 
    assign out[11084] = 1'b0; 
    assign out[11085] = 1'b0; 
    assign out[11086] = 1'b0; 
    assign out[11087] = 1'b0; 
    assign out[11088] = 1'b0; 
    assign out[11089] = 1'b0; 
    assign out[11090] = 1'b0; 
    assign out[11091] = 1'b0; 
    assign out[11092] = 1'b0; 
    assign out[11093] = 1'b0; 
    assign out[11094] = 1'b0; 
    assign out[11095] = 1'b0; 
    assign out[11096] = 1'b0; 
    assign out[11097] = 1'b0; 
    assign out[11098] = 1'b0; 
    assign out[11099] = 1'b0; 
    assign out[11100] = 1'b0; 
    assign out[11101] = 1'b0; 
    assign out[11102] = 1'b0; 
    assign out[11103] = 1'b0; 
    assign out[11104] = 1'b0; 
    assign out[11105] = 1'b0; 
    assign out[11106] = 1'b0; 
    assign out[11107] = 1'b0; 
    assign out[11108] = 1'b0; 
    assign out[11109] = 1'b0; 
    assign out[11110] = 1'b0; 
    assign out[11111] = 1'b0; 
    assign out[11112] = 1'b0; 
    assign out[11113] = 1'b0; 
    assign out[11114] = 1'b0; 
    assign out[11115] = 1'b0; 
    assign out[11116] = 1'b0; 
    assign out[11117] = 1'b0; 
    assign out[11118] = 1'b0; 
    assign out[11119] = 1'b0; 
    assign out[11120] = 1'b0; 
    assign out[11121] = 1'b0; 
    assign out[11122] = 1'b0; 
    assign out[11123] = 1'b0; 
    assign out[11124] = 1'b0; 
    assign out[11125] = 1'b0; 
    assign out[11126] = 1'b0; 
    assign out[11127] = 1'b0; 
    assign out[11128] = 1'b0; 
    assign out[11129] = 1'b0; 
    assign out[11130] = 1'b0; 
    assign out[11131] = 1'b0; 
    assign out[11132] = 1'b0; 
    assign out[11133] = 1'b0; 
    assign out[11134] = 1'b0; 
    assign out[11135] = 1'b0; 
    assign out[11136] = 1'b0; 
    assign out[11137] = 1'b0; 
    assign out[11138] = 1'b0; 
    assign out[11139] = 1'b0; 
    assign out[11140] = 1'b0; 
    assign out[11141] = 1'b0; 
    assign out[11142] = 1'b0; 
    assign out[11143] = 1'b0; 
    assign out[11144] = 1'b0; 
    assign out[11145] = 1'b0; 
    assign out[11146] = 1'b0; 
    assign out[11147] = 1'b0; 
    assign out[11148] = 1'b0; 
    assign out[11149] = 1'b0; 
    assign out[11150] = 1'b0; 
    assign out[11151] = 1'b0; 
    assign out[11152] = 1'b0; 
    assign out[11153] = 1'b0; 
    assign out[11154] = 1'b0; 
    assign out[11155] = 1'b0; 
    assign out[11156] = 1'b0; 
    assign out[11157] = 1'b0; 
    assign out[11158] = 1'b0; 
    assign out[11159] = 1'b0; 
    assign out[11160] = 1'b0; 
    assign out[11161] = 1'b0; 
    assign out[11162] = 1'b0; 
    assign out[11163] = 1'b0; 
    assign out[11164] = 1'b0; 
    assign out[11165] = 1'b0; 
    assign out[11166] = 1'b0; 
    assign out[11167] = 1'b0; 
    assign out[11168] = 1'b0; 
    assign out[11169] = 1'b0; 
    assign out[11170] = 1'b0; 
    assign out[11171] = 1'b0; 
    assign out[11172] = 1'b0; 
    assign out[11173] = 1'b0; 
    assign out[11174] = 1'b0; 
    assign out[11175] = 1'b0; 
    assign out[11176] = 1'b0; 
    assign out[11177] = 1'b0; 
    assign out[11178] = 1'b0; 
    assign out[11179] = 1'b0; 
    assign out[11180] = 1'b0; 
    assign out[11181] = 1'b0; 
    assign out[11182] = 1'b0; 
    assign out[11183] = 1'b0; 
    assign out[11184] = 1'b0; 
    assign out[11185] = 1'b0; 
    assign out[11186] = 1'b0; 
    assign out[11187] = 1'b0; 
    assign out[11188] = 1'b0; 
    assign out[11189] = 1'b0; 
    assign out[11190] = 1'b0; 
    assign out[11191] = 1'b0; 
    assign out[11192] = 1'b0; 
    assign out[11193] = 1'b0; 
    assign out[11194] = 1'b0; 
    assign out[11195] = 1'b0; 
    assign out[11196] = 1'b0; 
    assign out[11197] = 1'b0; 
    assign out[11198] = 1'b0; 
    assign out[11199] = 1'b0; 
    assign out[11200] = 1'b0; 
    assign out[11201] = 1'b0; 
    assign out[11202] = 1'b0; 
    assign out[11203] = 1'b0; 
    assign out[11204] = 1'b0; 
    assign out[11205] = 1'b0; 
    assign out[11206] = 1'b0; 
    assign out[11207] = 1'b0; 
    assign out[11208] = 1'b0; 
    assign out[11209] = 1'b0; 
    assign out[11210] = 1'b0; 
    assign out[11211] = 1'b0; 
    assign out[11212] = 1'b0; 
    assign out[11213] = 1'b0; 
    assign out[11214] = 1'b0; 
    assign out[11215] = 1'b0; 
    assign out[11216] = 1'b0; 
    assign out[11217] = 1'b0; 
    assign out[11218] = 1'b0; 
    assign out[11219] = 1'b0; 
    assign out[11220] = 1'b0; 
    assign out[11221] = 1'b0; 
    assign out[11222] = 1'b0; 
    assign out[11223] = 1'b0; 
    assign out[11224] = 1'b0; 
    assign out[11225] = 1'b0; 
    assign out[11226] = 1'b0; 
    assign out[11227] = 1'b0; 
    assign out[11228] = 1'b0; 
    assign out[11229] = 1'b0; 
    assign out[11230] = 1'b0; 
    assign out[11231] = 1'b0; 
    assign out[11232] = 1'b0; 
    assign out[11233] = 1'b0; 
    assign out[11234] = 1'b0; 
    assign out[11235] = 1'b0; 
    assign out[11236] = 1'b0; 
    assign out[11237] = 1'b0; 
    assign out[11238] = 1'b0; 
    assign out[11239] = 1'b0; 
    assign out[11240] = 1'b0; 
    assign out[11241] = 1'b0; 
    assign out[11242] = 1'b0; 
    assign out[11243] = 1'b0; 
    assign out[11244] = 1'b0; 
    assign out[11245] = 1'b0; 
    assign out[11246] = 1'b0; 
    assign out[11247] = 1'b0; 
    assign out[11248] = 1'b0; 
    assign out[11249] = 1'b0; 
    assign out[11250] = 1'b0; 
    assign out[11251] = 1'b0; 
    assign out[11252] = 1'b0; 
    assign out[11253] = 1'b0; 
    assign out[11254] = 1'b0; 
    assign out[11255] = 1'b0; 
    assign out[11256] = 1'b0; 
    assign out[11257] = 1'b0; 
    assign out[11258] = 1'b0; 
    assign out[11259] = 1'b0; 
    assign out[11260] = 1'b0; 
    assign out[11261] = 1'b0; 
    assign out[11262] = 1'b0; 
    assign out[11263] = 1'b0; 
    assign out[11264] = 1'b0; 
    assign out[11265] = 1'b0; 
    assign out[11266] = 1'b0; 
    assign out[11267] = 1'b0; 
    assign out[11268] = 1'b0; 
    assign out[11269] = 1'b0; 
    assign out[11270] = 1'b0; 
    assign out[11271] = 1'b0; 
    assign out[11272] = 1'b0; 
    assign out[11273] = 1'b0; 
    assign out[11274] = 1'b0; 
    assign out[11275] = 1'b0; 
    assign out[11276] = 1'b0; 
    assign out[11277] = 1'b0; 
    assign out[11278] = 1'b0; 
    assign out[11279] = 1'b0; 
    assign out[11280] = 1'b0; 
    assign out[11281] = 1'b0; 
    assign out[11282] = 1'b0; 
    assign out[11283] = 1'b0; 
    assign out[11284] = 1'b0; 
    assign out[11285] = 1'b0; 
    assign out[11286] = 1'b0; 
    assign out[11287] = 1'b0; 
    assign out[11288] = 1'b0; 
    assign out[11289] = 1'b0; 
    assign out[11290] = 1'b0; 
    assign out[11291] = 1'b0; 
    assign out[11292] = 1'b0; 
    assign out[11293] = 1'b0; 
    assign out[11294] = 1'b0; 
    assign out[11295] = 1'b0; 
    assign out[11296] = 1'b0; 
    assign out[11297] = 1'b0; 
    assign out[11298] = 1'b0; 
    assign out[11299] = 1'b0; 
    assign out[11300] = 1'b0; 
    assign out[11301] = 1'b0; 
    assign out[11302] = 1'b0; 
    assign out[11303] = 1'b0; 
    assign out[11304] = 1'b0; 
    assign out[11305] = 1'b0; 
    assign out[11306] = 1'b0; 
    assign out[11307] = 1'b0; 
    assign out[11308] = 1'b0; 
    assign out[11309] = 1'b0; 
    assign out[11310] = 1'b0; 
    assign out[11311] = 1'b0; 
    assign out[11312] = 1'b0; 
    assign out[11313] = 1'b0; 
    assign out[11314] = 1'b0; 
    assign out[11315] = 1'b0; 
    assign out[11316] = 1'b0; 
    assign out[11317] = 1'b0; 
    assign out[11318] = 1'b0; 
    assign out[11319] = 1'b0; 
    assign out[11320] = 1'b0; 
    assign out[11321] = 1'b0; 
    assign out[11322] = 1'b0; 
    assign out[11323] = 1'b0; 
    assign out[11324] = 1'b0; 
    assign out[11325] = 1'b0; 
    assign out[11326] = 1'b0; 
    assign out[11327] = 1'b0; 
    assign out[11328] = 1'b0; 
    assign out[11329] = 1'b0; 
    assign out[11330] = 1'b0; 
    assign out[11331] = 1'b0; 
    assign out[11332] = 1'b0; 
    assign out[11333] = 1'b0; 
    assign out[11334] = 1'b0; 
    assign out[11335] = 1'b0; 
    assign out[11336] = 1'b0; 
    assign out[11337] = 1'b0; 
    assign out[11338] = 1'b0; 
    assign out[11339] = 1'b0; 
    assign out[11340] = 1'b0; 
    assign out[11341] = 1'b0; 
    assign out[11342] = 1'b0; 
    assign out[11343] = 1'b0; 
    assign out[11344] = 1'b0; 
    assign out[11345] = 1'b0; 
    assign out[11346] = 1'b0; 
    assign out[11347] = 1'b0; 
    assign out[11348] = 1'b0; 
    assign out[11349] = 1'b0; 
    assign out[11350] = 1'b0; 
    assign out[11351] = 1'b0; 
    assign out[11352] = 1'b0; 
    assign out[11353] = 1'b0; 
    assign out[11354] = 1'b0; 
    assign out[11355] = 1'b0; 
    assign out[11356] = 1'b0; 
    assign out[11357] = 1'b0; 
    assign out[11358] = 1'b0; 
    assign out[11359] = 1'b0; 
    assign out[11360] = 1'b0; 
    assign out[11361] = 1'b0; 
    assign out[11362] = 1'b0; 
    assign out[11363] = 1'b0; 
    assign out[11364] = 1'b0; 
    assign out[11365] = 1'b0; 
    assign out[11366] = 1'b0; 
    assign out[11367] = 1'b0; 
    assign out[11368] = 1'b0; 
    assign out[11369] = 1'b0; 
    assign out[11370] = 1'b0; 
    assign out[11371] = 1'b0; 
    assign out[11372] = 1'b0; 
    assign out[11373] = 1'b0; 
    assign out[11374] = 1'b0; 
    assign out[11375] = 1'b0; 
    assign out[11376] = 1'b0; 
    assign out[11377] = 1'b0; 
    assign out[11378] = 1'b0; 
    assign out[11379] = 1'b0; 
    assign out[11380] = 1'b0; 
    assign out[11381] = 1'b0; 
    assign out[11382] = 1'b0; 
    assign out[11383] = 1'b0; 
    assign out[11384] = 1'b0; 
    assign out[11385] = 1'b0; 
    assign out[11386] = 1'b0; 
    assign out[11387] = 1'b0; 
    assign out[11388] = 1'b0; 
    assign out[11389] = 1'b0; 
    assign out[11390] = 1'b0; 
    assign out[11391] = 1'b0; 
    assign out[11392] = 1'b0; 
    assign out[11393] = 1'b0; 
    assign out[11394] = 1'b0; 
    assign out[11395] = 1'b0; 
    assign out[11396] = 1'b0; 
    assign out[11397] = 1'b0; 
    assign out[11398] = 1'b0; 
    assign out[11399] = 1'b0; 
    assign out[11400] = 1'b0; 
    assign out[11401] = 1'b0; 
    assign out[11402] = 1'b0; 
    assign out[11403] = 1'b0; 
    assign out[11404] = 1'b0; 
    assign out[11405] = 1'b0; 
    assign out[11406] = 1'b0; 
    assign out[11407] = 1'b0; 
    assign out[11408] = 1'b0; 
    assign out[11409] = 1'b0; 
    assign out[11410] = 1'b0; 
    assign out[11411] = 1'b0; 
    assign out[11412] = 1'b0; 
    assign out[11413] = 1'b0; 
    assign out[11414] = 1'b0; 
    assign out[11415] = 1'b0; 
    assign out[11416] = 1'b0; 
    assign out[11417] = 1'b0; 
    assign out[11418] = 1'b0; 
    assign out[11419] = 1'b0; 
    assign out[11420] = 1'b0; 
    assign out[11421] = 1'b0; 
    assign out[11422] = 1'b0; 
    assign out[11423] = 1'b0; 
    assign out[11424] = 1'b0; 
    assign out[11425] = 1'b0; 
    assign out[11426] = 1'b0; 
    assign out[11427] = 1'b0; 
    assign out[11428] = 1'b0; 
    assign out[11429] = 1'b0; 
    assign out[11430] = 1'b0; 
    assign out[11431] = 1'b0; 
    assign out[11432] = 1'b0; 
    assign out[11433] = 1'b0; 
    assign out[11434] = 1'b0; 
    assign out[11435] = 1'b0; 
    assign out[11436] = 1'b0; 
    assign out[11437] = 1'b0; 
    assign out[11438] = 1'b0; 
    assign out[11439] = 1'b0; 
    assign out[11440] = 1'b0; 
    assign out[11441] = 1'b0; 
    assign out[11442] = 1'b0; 
    assign out[11443] = 1'b0; 
    assign out[11444] = 1'b0; 
    assign out[11445] = 1'b0; 
    assign out[11446] = 1'b0; 
    assign out[11447] = 1'b0; 
    assign out[11448] = 1'b0; 
    assign out[11449] = 1'b0; 
    assign out[11450] = 1'b0; 
    assign out[11451] = 1'b0; 
    assign out[11452] = 1'b0; 
    assign out[11453] = 1'b0; 
    assign out[11454] = 1'b0; 
    assign out[11455] = 1'b0; 
    assign out[11456] = 1'b0; 
    assign out[11457] = 1'b0; 
    assign out[11458] = 1'b0; 
    assign out[11459] = 1'b0; 
    assign out[11460] = 1'b0; 
    assign out[11461] = 1'b0; 
    assign out[11462] = 1'b0; 
    assign out[11463] = 1'b0; 
    assign out[11464] = 1'b0; 
    assign out[11465] = 1'b0; 
    assign out[11466] = 1'b0; 
    assign out[11467] = 1'b0; 
    assign out[11468] = 1'b0; 
    assign out[11469] = 1'b0; 
    assign out[11470] = 1'b0; 
    assign out[11471] = 1'b0; 
    assign out[11472] = 1'b0; 
    assign out[11473] = 1'b0; 
    assign out[11474] = 1'b0; 
    assign out[11475] = 1'b0; 
    assign out[11476] = 1'b0; 
    assign out[11477] = 1'b0; 
    assign out[11478] = 1'b0; 
    assign out[11479] = 1'b0; 
    assign out[11480] = 1'b0; 
    assign out[11481] = 1'b0; 
    assign out[11482] = 1'b0; 
    assign out[11483] = 1'b0; 
    assign out[11484] = 1'b0; 
    assign out[11485] = 1'b0; 
    assign out[11486] = 1'b0; 
    assign out[11487] = 1'b0; 
    assign out[11488] = 1'b0; 
    assign out[11489] = 1'b0; 
    assign out[11490] = 1'b0; 
    assign out[11491] = 1'b0; 
    assign out[11492] = 1'b0; 
    assign out[11493] = 1'b0; 
    assign out[11494] = 1'b0; 
    assign out[11495] = 1'b0; 
    assign out[11496] = 1'b0; 
    assign out[11497] = 1'b0; 
    assign out[11498] = 1'b0; 
    assign out[11499] = 1'b0; 
    assign out[11500] = 1'b0; 
    assign out[11501] = 1'b0; 
    assign out[11502] = 1'b0; 
    assign out[11503] = 1'b0; 
    assign out[11504] = 1'b0; 
    assign out[11505] = 1'b0; 
    assign out[11506] = 1'b0; 
    assign out[11507] = 1'b0; 
    assign out[11508] = 1'b0; 
    assign out[11509] = 1'b0; 
    assign out[11510] = 1'b0; 
    assign out[11511] = 1'b0; 
    assign out[11512] = 1'b0; 
    assign out[11513] = 1'b0; 
    assign out[11514] = 1'b0; 
    assign out[11515] = 1'b0; 
    assign out[11516] = 1'b0; 
    assign out[11517] = 1'b0; 
    assign out[11518] = 1'b0; 
    assign out[11519] = 1'b0; 
    assign out[11520] = 1'b0; 
    assign out[11521] = 1'b0; 
    assign out[11522] = 1'b0; 
    assign out[11523] = 1'b0; 
    assign out[11524] = 1'b0; 
    assign out[11525] = 1'b0; 
    assign out[11526] = 1'b0; 
    assign out[11527] = 1'b0; 
    assign out[11528] = 1'b0; 
    assign out[11529] = 1'b0; 
    assign out[11530] = 1'b0; 
    assign out[11531] = 1'b0; 
    assign out[11532] = 1'b0; 
    assign out[11533] = 1'b0; 
    assign out[11534] = 1'b0; 
    assign out[11535] = 1'b0; 
    assign out[11536] = 1'b0; 
    assign out[11537] = 1'b0; 
    assign out[11538] = 1'b0; 
    assign out[11539] = 1'b0; 
    assign out[11540] = 1'b0; 
    assign out[11541] = 1'b0; 
    assign out[11542] = 1'b0; 
    assign out[11543] = 1'b0; 
    assign out[11544] = 1'b0; 
    assign out[11545] = 1'b0; 
    assign out[11546] = 1'b0; 
    assign out[11547] = 1'b0; 
    assign out[11548] = 1'b0; 
    assign out[11549] = 1'b0; 
    assign out[11550] = 1'b0; 
    assign out[11551] = 1'b0; 
    assign out[11552] = 1'b0; 
    assign out[11553] = 1'b0; 
    assign out[11554] = 1'b0; 
    assign out[11555] = 1'b0; 
    assign out[11556] = 1'b0; 
    assign out[11557] = 1'b0; 
    assign out[11558] = 1'b0; 
    assign out[11559] = 1'b0; 
    assign out[11560] = 1'b0; 
    assign out[11561] = 1'b0; 
    assign out[11562] = 1'b0; 
    assign out[11563] = 1'b0; 
    assign out[11564] = 1'b0; 
    assign out[11565] = 1'b0; 
    assign out[11566] = 1'b0; 
    assign out[11567] = 1'b0; 
    assign out[11568] = 1'b0; 
    assign out[11569] = 1'b0; 
    assign out[11570] = 1'b0; 
    assign out[11571] = 1'b0; 
    assign out[11572] = 1'b0; 
    assign out[11573] = 1'b0; 
    assign out[11574] = 1'b0; 
    assign out[11575] = 1'b0; 
    assign out[11576] = 1'b0; 
    assign out[11577] = 1'b0; 
    assign out[11578] = 1'b0; 
    assign out[11579] = 1'b0; 
    assign out[11580] = 1'b0; 
    assign out[11581] = 1'b0; 
    assign out[11582] = 1'b0; 
    assign out[11583] = 1'b0; 
    assign out[11584] = 1'b0; 
    assign out[11585] = 1'b0; 
    assign out[11586] = 1'b0; 
    assign out[11587] = 1'b0; 
    assign out[11588] = 1'b0; 
    assign out[11589] = 1'b0; 
    assign out[11590] = 1'b0; 
    assign out[11591] = 1'b0; 
    assign out[11592] = 1'b0; 
    assign out[11593] = 1'b0; 
    assign out[11594] = 1'b0; 
    assign out[11595] = 1'b0; 
    assign out[11596] = 1'b0; 
    assign out[11597] = 1'b0; 
    assign out[11598] = 1'b0; 
    assign out[11599] = 1'b0; 
    assign out[11600] = 1'b0; 
    assign out[11601] = 1'b0; 
    assign out[11602] = 1'b0; 
    assign out[11603] = 1'b0; 
    assign out[11604] = 1'b0; 
    assign out[11605] = 1'b0; 
    assign out[11606] = 1'b0; 
    assign out[11607] = 1'b0; 
    assign out[11608] = 1'b0; 
    assign out[11609] = 1'b0; 
    assign out[11610] = 1'b0; 
    assign out[11611] = 1'b0; 
    assign out[11612] = 1'b0; 
    assign out[11613] = 1'b0; 
    assign out[11614] = 1'b0; 
    assign out[11615] = 1'b0; 
    assign out[11616] = 1'b0; 
    assign out[11617] = 1'b0; 
    assign out[11618] = 1'b0; 
    assign out[11619] = 1'b0; 
    assign out[11620] = 1'b0; 
    assign out[11621] = 1'b0; 
    assign out[11622] = 1'b0; 
    assign out[11623] = 1'b0; 
    assign out[11624] = 1'b0; 
    assign out[11625] = 1'b0; 
    assign out[11626] = 1'b0; 
    assign out[11627] = 1'b0; 
    assign out[11628] = 1'b0; 
    assign out[11629] = 1'b0; 
    assign out[11630] = 1'b0; 
    assign out[11631] = 1'b0; 
    assign out[11632] = 1'b0; 
    assign out[11633] = 1'b0; 
    assign out[11634] = 1'b0; 
    assign out[11635] = 1'b0; 
    assign out[11636] = 1'b0; 
    assign out[11637] = 1'b0; 
    assign out[11638] = 1'b0; 
    assign out[11639] = 1'b0; 
    assign out[11640] = 1'b0; 
    assign out[11641] = 1'b0; 
    assign out[11642] = 1'b0; 
    assign out[11643] = 1'b0; 
    assign out[11644] = 1'b0; 
    assign out[11645] = 1'b0; 
    assign out[11646] = 1'b0; 
    assign out[11647] = 1'b0; 
    assign out[11648] = 1'b0; 
    assign out[11649] = 1'b0; 
    assign out[11650] = 1'b0; 
    assign out[11651] = 1'b0; 
    assign out[11652] = 1'b0; 
    assign out[11653] = 1'b0; 
    assign out[11654] = 1'b0; 
    assign out[11655] = 1'b0; 
    assign out[11656] = 1'b0; 
    assign out[11657] = 1'b0; 
    assign out[11658] = 1'b0; 
    assign out[11659] = 1'b0; 
    assign out[11660] = 1'b0; 
    assign out[11661] = 1'b0; 
    assign out[11662] = 1'b0; 
    assign out[11663] = 1'b0; 
    assign out[11664] = 1'b0; 
    assign out[11665] = 1'b0; 
    assign out[11666] = 1'b0; 
    assign out[11667] = 1'b0; 
    assign out[11668] = 1'b0; 
    assign out[11669] = 1'b0; 
    assign out[11670] = 1'b0; 
    assign out[11671] = 1'b0; 
    assign out[11672] = 1'b0; 
    assign out[11673] = 1'b0; 
    assign out[11674] = 1'b0; 
    assign out[11675] = 1'b0; 
    assign out[11676] = 1'b0; 
    assign out[11677] = 1'b0; 
    assign out[11678] = 1'b0; 
    assign out[11679] = 1'b0; 
    assign out[11680] = 1'b0; 
    assign out[11681] = 1'b0; 
    assign out[11682] = 1'b0; 
    assign out[11683] = 1'b0; 
    assign out[11684] = 1'b0; 
    assign out[11685] = 1'b0; 
    assign out[11686] = 1'b0; 
    assign out[11687] = 1'b0; 
    assign out[11688] = 1'b0; 
    assign out[11689] = 1'b0; 
    assign out[11690] = 1'b0; 
    assign out[11691] = 1'b0; 
    assign out[11692] = 1'b0; 
    assign out[11693] = 1'b0; 
    assign out[11694] = 1'b0; 
    assign out[11695] = 1'b0; 
    assign out[11696] = 1'b0; 
    assign out[11697] = 1'b0; 
    assign out[11698] = 1'b0; 
    assign out[11699] = 1'b0; 
    assign out[11700] = 1'b0; 
    assign out[11701] = 1'b0; 
    assign out[11702] = 1'b0; 
    assign out[11703] = 1'b0; 
    assign out[11704] = 1'b0; 
    assign out[11705] = 1'b0; 
    assign out[11706] = 1'b0; 
    assign out[11707] = 1'b0; 
    assign out[11708] = 1'b0; 
    assign out[11709] = 1'b0; 
    assign out[11710] = 1'b0; 
    assign out[11711] = 1'b0; 
    assign out[11712] = 1'b0; 
    assign out[11713] = 1'b0; 
    assign out[11714] = 1'b0; 
    assign out[11715] = 1'b0; 
    assign out[11716] = 1'b0; 
    assign out[11717] = 1'b0; 
    assign out[11718] = 1'b0; 
    assign out[11719] = 1'b0; 
    assign out[11720] = 1'b0; 
    assign out[11721] = 1'b0; 
    assign out[11722] = 1'b0; 
    assign out[11723] = 1'b0; 
    assign out[11724] = 1'b0; 
    assign out[11725] = 1'b0; 
    assign out[11726] = 1'b0; 
    assign out[11727] = 1'b0; 
    assign out[11728] = 1'b0; 
    assign out[11729] = 1'b0; 
    assign out[11730] = 1'b0; 
    assign out[11731] = 1'b0; 
    assign out[11732] = 1'b0; 
    assign out[11733] = 1'b0; 
    assign out[11734] = 1'b0; 
    assign out[11735] = 1'b0; 
    assign out[11736] = 1'b0; 
    assign out[11737] = 1'b0; 
    assign out[11738] = 1'b0; 
    assign out[11739] = 1'b0; 
    assign out[11740] = 1'b0; 
    assign out[11741] = 1'b0; 
    assign out[11742] = 1'b0; 
    assign out[11743] = 1'b0; 
    assign out[11744] = 1'b0; 
    assign out[11745] = 1'b0; 
    assign out[11746] = 1'b0; 
    assign out[11747] = 1'b0; 
    assign out[11748] = 1'b0; 
    assign out[11749] = 1'b0; 
    assign out[11750] = 1'b0; 
    assign out[11751] = 1'b0; 
    assign out[11752] = 1'b0; 
    assign out[11753] = 1'b0; 
    assign out[11754] = 1'b0; 
    assign out[11755] = 1'b0; 
    assign out[11756] = 1'b0; 
    assign out[11757] = 1'b0; 
    assign out[11758] = 1'b0; 
    assign out[11759] = 1'b0; 
    assign out[11760] = 1'b0; 
    assign out[11761] = 1'b0; 
    assign out[11762] = 1'b0; 
    assign out[11763] = 1'b0; 
    assign out[11764] = 1'b0; 
    assign out[11765] = 1'b0; 
    assign out[11766] = 1'b0; 
    assign out[11767] = 1'b0; 
    assign out[11768] = 1'b0; 
    assign out[11769] = 1'b0; 
    assign out[11770] = 1'b0; 
    assign out[11771] = 1'b0; 
    assign out[11772] = 1'b0; 
    assign out[11773] = 1'b0; 
    assign out[11774] = 1'b0; 
    assign out[11775] = 1'b0; 
    assign out[11776] = 1'b0; 
    assign out[11777] = 1'b0; 
    assign out[11778] = 1'b0; 
    assign out[11779] = 1'b0; 
    assign out[11780] = 1'b0; 
    assign out[11781] = 1'b0; 
    assign out[11782] = 1'b0; 
    assign out[11783] = 1'b0; 
    assign out[11784] = 1'b0; 
    assign out[11785] = 1'b0; 
    assign out[11786] = 1'b0; 
    assign out[11787] = 1'b0; 
    assign out[11788] = 1'b0; 
    assign out[11789] = 1'b0; 
    assign out[11790] = 1'b0; 
    assign out[11791] = 1'b0; 
    assign out[11792] = 1'b0; 
    assign out[11793] = 1'b0; 
    assign out[11794] = 1'b0; 
    assign out[11795] = 1'b0; 
    assign out[11796] = 1'b0; 
    assign out[11797] = 1'b0; 
    assign out[11798] = 1'b0; 
    assign out[11799] = 1'b0; 
    assign out[11800] = 1'b0; 
    assign out[11801] = 1'b0; 
    assign out[11802] = 1'b0; 
    assign out[11803] = 1'b0; 
    assign out[11804] = 1'b0; 
    assign out[11805] = 1'b0; 
    assign out[11806] = 1'b0; 
    assign out[11807] = 1'b0; 
    assign out[11808] = 1'b0; 
    assign out[11809] = 1'b0; 
    assign out[11810] = 1'b0; 
    assign out[11811] = 1'b0; 
    assign out[11812] = 1'b0; 
    assign out[11813] = 1'b0; 
    assign out[11814] = 1'b0; 
    assign out[11815] = 1'b0; 
    assign out[11816] = 1'b0; 
    assign out[11817] = 1'b0; 
    assign out[11818] = 1'b0; 
    assign out[11819] = 1'b0; 
    assign out[11820] = 1'b0; 
    assign out[11821] = 1'b0; 
    assign out[11822] = 1'b0; 
    assign out[11823] = 1'b0; 
    assign out[11824] = 1'b0; 
    assign out[11825] = 1'b0; 
    assign out[11826] = 1'b0; 
    assign out[11827] = 1'b0; 
    assign out[11828] = 1'b0; 
    assign out[11829] = 1'b0; 
    assign out[11830] = 1'b0; 
    assign out[11831] = 1'b0; 
    assign out[11832] = 1'b0; 
    assign out[11833] = 1'b0; 
    assign out[11834] = 1'b0; 
    assign out[11835] = 1'b0; 
    assign out[11836] = 1'b0; 
    assign out[11837] = 1'b0; 
    assign out[11838] = 1'b0; 
    assign out[11839] = 1'b0; 
    assign out[11840] = 1'b0; 
    assign out[11841] = 1'b0; 
    assign out[11842] = 1'b0; 
    assign out[11843] = 1'b0; 
    assign out[11844] = 1'b0; 
    assign out[11845] = 1'b0; 
    assign out[11846] = 1'b0; 
    assign out[11847] = 1'b0; 
    assign out[11848] = 1'b0; 
    assign out[11849] = 1'b0; 
    assign out[11850] = 1'b0; 
    assign out[11851] = 1'b0; 
    assign out[11852] = 1'b0; 
    assign out[11853] = 1'b0; 
    assign out[11854] = 1'b0; 
    assign out[11855] = 1'b0; 
    assign out[11856] = 1'b0; 
    assign out[11857] = 1'b0; 
    assign out[11858] = 1'b0; 
    assign out[11859] = 1'b0; 
    assign out[11860] = 1'b0; 
    assign out[11861] = 1'b0; 
    assign out[11862] = 1'b0; 
    assign out[11863] = 1'b0; 
    assign out[11864] = 1'b0; 
    assign out[11865] = 1'b0; 
    assign out[11866] = 1'b0; 
    assign out[11867] = 1'b0; 
    assign out[11868] = 1'b0; 
    assign out[11869] = 1'b0; 
    assign out[11870] = 1'b0; 
    assign out[11871] = 1'b0; 
    assign out[11872] = 1'b0; 
    assign out[11873] = 1'b0; 
    assign out[11874] = 1'b0; 
    assign out[11875] = 1'b0; 
    assign out[11876] = 1'b0; 
    assign out[11877] = 1'b0; 
    assign out[11878] = 1'b0; 
    assign out[11879] = 1'b0; 
    assign out[11880] = 1'b0; 
    assign out[11881] = 1'b0; 
    assign out[11882] = 1'b0; 
    assign out[11883] = 1'b0; 
    assign out[11884] = 1'b0; 
    assign out[11885] = 1'b0; 
    assign out[11886] = 1'b0; 
    assign out[11887] = 1'b0; 
    assign out[11888] = 1'b0; 
    assign out[11889] = 1'b0; 
    assign out[11890] = 1'b0; 
    assign out[11891] = 1'b0; 
    assign out[11892] = 1'b0; 
    assign out[11893] = 1'b0; 
    assign out[11894] = 1'b0; 
    assign out[11895] = 1'b0; 
    assign out[11896] = 1'b0; 
    assign out[11897] = 1'b0; 
    assign out[11898] = 1'b0; 
    assign out[11899] = 1'b0; 
    assign out[11900] = 1'b0; 
    assign out[11901] = 1'b0; 
    assign out[11902] = 1'b0; 
    assign out[11903] = 1'b0; 
    assign out[11904] = 1'b0; 
    assign out[11905] = 1'b0; 
    assign out[11906] = 1'b0; 
    assign out[11907] = 1'b0; 
    assign out[11908] = 1'b0; 
    assign out[11909] = 1'b0; 
    assign out[11910] = 1'b0; 
    assign out[11911] = 1'b0; 
    assign out[11912] = 1'b0; 
    assign out[11913] = 1'b0; 
    assign out[11914] = 1'b0; 
    assign out[11915] = 1'b0; 
    assign out[11916] = 1'b0; 
    assign out[11917] = 1'b0; 
    assign out[11918] = 1'b0; 
    assign out[11919] = 1'b0; 
    assign out[11920] = 1'b0; 
    assign out[11921] = 1'b0; 
    assign out[11922] = 1'b0; 
    assign out[11923] = 1'b0; 
    assign out[11924] = 1'b0; 
    assign out[11925] = 1'b0; 
    assign out[11926] = 1'b0; 
    assign out[11927] = 1'b0; 
    assign out[11928] = 1'b0; 
    assign out[11929] = 1'b0; 
    assign out[11930] = 1'b0; 
    assign out[11931] = 1'b0; 
    assign out[11932] = 1'b0; 
    assign out[11933] = 1'b0; 
    assign out[11934] = 1'b0; 
    assign out[11935] = 1'b0; 
    assign out[11936] = 1'b0; 
    assign out[11937] = 1'b0; 
    assign out[11938] = 1'b0; 
    assign out[11939] = 1'b0; 
    assign out[11940] = 1'b0; 
    assign out[11941] = 1'b0; 
    assign out[11942] = 1'b0; 
    assign out[11943] = 1'b0; 
    assign out[11944] = 1'b0; 
    assign out[11945] = 1'b0; 
    assign out[11946] = 1'b0; 
    assign out[11947] = 1'b0; 
    assign out[11948] = 1'b0; 
    assign out[11949] = 1'b0; 
    assign out[11950] = 1'b0; 
    assign out[11951] = 1'b0; 
    assign out[11952] = 1'b0; 
    assign out[11953] = 1'b0; 
    assign out[11954] = 1'b0; 
    assign out[11955] = 1'b0; 
    assign out[11956] = 1'b0; 
    assign out[11957] = 1'b0; 
    assign out[11958] = 1'b0; 
    assign out[11959] = 1'b0; 
    assign out[11960] = 1'b0; 
    assign out[11961] = 1'b0; 
    assign out[11962] = 1'b0; 
    assign out[11963] = 1'b0; 
    assign out[11964] = 1'b0; 
    assign out[11965] = 1'b0; 
    assign out[11966] = 1'b0; 
    assign out[11967] = 1'b0; 
    assign out[11968] = 1'b0; 
    assign out[11969] = 1'b0; 
    assign out[11970] = 1'b0; 
    assign out[11971] = 1'b0; 
    assign out[11972] = 1'b0; 
    assign out[11973] = 1'b0; 
    assign out[11974] = 1'b0; 
    assign out[11975] = 1'b0; 
    assign out[11976] = 1'b0; 
    assign out[11977] = 1'b0; 
    assign out[11978] = 1'b0; 
    assign out[11979] = 1'b0; 
    assign out[11980] = 1'b0; 
    assign out[11981] = 1'b0; 
    assign out[11982] = 1'b0; 
    assign out[11983] = 1'b0; 
    assign out[11984] = 1'b0; 
    assign out[11985] = 1'b0; 
    assign out[11986] = 1'b0; 
    assign out[11987] = 1'b0; 
    assign out[11988] = 1'b0; 
    assign out[11989] = 1'b0; 
    assign out[11990] = 1'b0; 
    assign out[11991] = 1'b0; 
    assign out[11992] = 1'b0; 
    assign out[11993] = 1'b0; 
    assign out[11994] = 1'b0; 
    assign out[11995] = 1'b0; 
    assign out[11996] = 1'b0; 
    assign out[11997] = 1'b0; 
    assign out[11998] = 1'b0; 
    assign out[11999] = 1'b0; 
    // Arrange outputs in categories ================================================
    assign categories[7999:0] = out[7999:0];

endmodule
